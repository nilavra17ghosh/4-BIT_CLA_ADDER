* SPICE3 file created from xor1.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale=0.09u
.global gnd vdd

VDS vdd gnd 'SUPPLY'
vin1 A gnd pulse 0 1.8 0ns 100ps 100ps 9.9ns 20ns
vin2 B gnd pulse 0 1.8 0ns 100ps 100ps 19.9ns 40ns

M1000 a_24_2# B XOR VDD CMOSP w=6 l=2
+  ad=48 pd=28 as=48 ps=28
M1001 VDD A Anot VDD CMOSP w=6 l=2
+  ad=120 pd=88 as=30 ps=22
M1002 GND A Anot Gnd CMOSN w=4 l=2
+  ad=80 pd=72 as=20 ps=18
M1003 XOR Bnot a_4_2# VDD CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1004 Bnot B GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 GND Anot a_24_n44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1006 a_4_2# A VDD VDD CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_24_n44# Bnot XOR Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1008 VDD Anot a_24_2# VDD CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 XOR B a_4_n44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1010 a_4_n44# A GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 Bnot B VDD VDD CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0

C0 XOR B 0.01fF
C1 B VDD 0.23fF
C2 B GND 0.08fF
C3 B Bnot 0.08fF
C4 A VDD 0.13fF
C5 XOR VDD 0.02fF
C6 VDD VDD 0.12fF
C7 B Anot 0.10fF
C8 XOR A 0.10fF
C9 Bnot VDD 0.09fF
C10 A GND 0.12fF
C11 A Bnot 0.20fF
C12 XOR Bnot 0.12fF
C13 Bnot VDD 0.12fF
C14 Anot VDD 0.09fF
C15 Bnot GND 0.08fF
C16 A Anot 0.28fF
C17 XOR Anot 0.09fF
C18 Anot VDD 0.06fF
C19 Anot GND 0.04fF
C20 B VDD 0.14fF
C21 B A 0.64fF
C22 GND Gnd 0.45fF
C23 XOR Gnd 0.58fF
C24 VDD Gnd 0.36fF
C25 Anot Gnd 0.42fF
C26 Bnot Gnd 0.50fF
C27 A Gnd 1.71fF
C28 B Gnd 1.24fF
C29 VDD Gnd 1.63fF

.tran 0.01n 80n

.control
run

set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
plot (v(XOR)+4) (v(A)+2) (v(B))

.endc
