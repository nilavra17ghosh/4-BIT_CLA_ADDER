magic
tech scmos
timestamp 1638596374
<< nwell >>
rect 0 -1 55 17
rect 61 -1 85 17
<< ntransistor >>
rect 11 -36 13 -32
rect 21 -36 23 -32
rect 31 -36 33 -32
rect 41 -36 43 -32
rect 72 -36 74 -32
<< ptransistor >>
rect 11 5 13 11
rect 21 5 23 11
rect 31 5 33 11
rect 41 5 43 11
rect 72 5 74 11
<< ndiffusion >>
rect 10 -36 11 -32
rect 13 -36 21 -32
rect 23 -36 31 -32
rect 33 -36 41 -32
rect 43 -36 45 -32
rect 71 -36 72 -32
rect 74 -36 75 -32
<< pdiffusion >>
rect 10 5 11 11
rect 13 5 15 11
rect 19 5 21 11
rect 23 5 25 11
rect 29 5 31 11
rect 33 5 35 11
rect 39 5 41 11
rect 43 5 45 11
rect 71 5 72 11
rect 74 5 75 11
<< ndcontact >>
rect 6 -36 10 -32
rect 45 -36 49 -32
rect 67 -36 71 -32
rect 75 -36 79 -32
<< pdcontact >>
rect 6 5 10 11
rect 15 5 19 11
rect 25 5 29 11
rect 35 5 39 11
rect 45 5 49 11
rect 67 5 71 11
rect 75 5 79 11
<< polysilicon >>
rect 11 11 13 20
rect 21 11 23 20
rect 31 11 33 20
rect 41 11 43 20
rect 72 11 74 20
rect 11 -32 13 5
rect 21 -32 23 5
rect 31 -32 33 5
rect 41 -32 43 5
rect 72 -32 74 5
rect 11 -39 13 -36
rect 21 -39 23 -36
rect 31 -39 33 -36
rect 41 -39 43 -36
rect 72 -39 74 -36
<< polycontact >>
rect 7 -7 11 -3
rect 17 -14 21 -10
rect 27 -21 31 -17
rect 37 -28 41 -24
rect 68 -7 72 -3
<< metal1 >>
rect 0 26 85 30
rect 6 11 10 26
rect 25 11 29 26
rect 45 11 49 26
rect 67 11 71 26
rect 15 -3 19 5
rect 35 -3 39 5
rect 75 -3 79 5
rect -5 -7 7 -3
rect 15 -7 68 -3
rect 75 -7 89 -3
rect -5 -14 17 -10
rect -5 -21 27 -17
rect -5 -28 37 -24
rect 45 -32 49 -7
rect 75 -32 79 -7
rect 6 -43 10 -36
rect 67 -43 71 -36
rect -1 -47 86 -43
<< end >>
