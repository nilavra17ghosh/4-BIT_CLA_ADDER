magic
tech scmos
timestamp 1637099764
<< nwell >>
rect 0 -1 37 17
rect 43 -1 67 17
<< ntransistor >>
rect 11 -25 13 -21
rect 21 -25 23 -21
rect 54 -25 56 -21
<< ptransistor >>
rect 11 5 13 11
rect 21 5 23 11
rect 54 5 56 11
<< ndiffusion >>
rect 10 -25 11 -21
rect 13 -25 21 -21
rect 23 -25 25 -21
rect 53 -25 54 -21
rect 56 -25 57 -21
<< pdiffusion >>
rect 10 5 11 11
rect 13 5 15 11
rect 19 5 21 11
rect 23 5 25 11
rect 53 5 54 11
rect 56 5 57 11
<< ndcontact >>
rect 6 -25 10 -21
rect 25 -25 29 -21
rect 49 -25 53 -21
rect 57 -25 61 -21
<< pdcontact >>
rect 6 5 10 11
rect 15 5 19 11
rect 25 5 29 11
rect 49 5 53 11
rect 57 5 61 11
<< polysilicon >>
rect 11 11 13 20
rect 21 11 23 20
rect 54 11 56 20
rect 11 -21 13 5
rect 21 -21 23 5
rect 54 -21 56 5
rect 11 -28 13 -25
rect 21 -28 23 -25
rect 54 -28 56 -25
<< polycontact >>
rect 7 -7 11 -3
rect 17 -16 21 -12
rect 50 -7 54 -3
<< metal1 >>
rect 0 26 67 29
rect 6 11 10 26
rect 25 11 29 26
rect 49 11 53 26
rect 15 -3 19 5
rect 57 -3 61 5
rect -5 -7 7 -3
rect 15 -7 50 -3
rect 57 -7 71 -3
rect -5 -16 17 -12
rect 25 -21 29 -7
rect 57 -21 61 -7
rect 6 -32 10 -25
rect 49 -32 53 -25
rect -1 -35 68 -32
<< labels >>
rlabel metal1 -5 -16 21 -12 1 B
rlabel metal1 -5 -7 11 -3 1 A
rlabel metal1 57 -7 71 -3 1 OUT
rlabel metal1 0 26 67 29 5 VDD
rlabel metal1 -1 -35 68 -32 1 GND
<< end >>
