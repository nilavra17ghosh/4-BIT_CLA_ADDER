magic
tech scmos
timestamp 1638569441
<< nwell >>
rect -13 7 73 25
<< ntransistor >>
rect -2 -44 0 -40
rect 8 -44 10 -40
rect 17 -44 19 -40
rect 27 -44 29 -40
rect 37 -44 39 -40
rect 55 -44 57 -40
<< ptransistor >>
rect -2 13 0 19
rect 8 13 10 19
rect 17 13 19 19
rect 27 13 29 19
rect 37 13 39 19
rect 55 13 57 19
<< ndiffusion >>
rect -3 -44 -2 -40
rect 0 -44 2 -40
rect 6 -44 8 -40
rect 10 -44 11 -40
rect 15 -44 17 -40
rect 19 -44 21 -40
rect 25 -44 27 -40
rect 29 -44 31 -40
rect 35 -44 37 -40
rect 39 -44 41 -40
rect 54 -44 55 -40
rect 57 -44 58 -40
<< pdiffusion >>
rect -3 13 -2 19
rect 0 13 8 19
rect 10 13 17 19
rect 19 13 27 19
rect 29 13 37 19
rect 39 13 41 19
rect 54 13 55 19
rect 57 13 58 19
<< ndcontact >>
rect -7 -44 -3 -40
rect 2 -44 6 -40
rect 11 -44 15 -40
rect 21 -44 25 -40
rect 31 -44 35 -40
rect 41 -44 45 -40
rect 50 -44 54 -40
rect 58 -44 62 -40
<< pdcontact >>
rect -7 13 -3 19
rect 41 13 45 19
rect 50 13 54 19
rect 58 13 62 19
<< polysilicon >>
rect -2 19 0 22
rect 8 19 10 22
rect 17 19 19 22
rect 27 19 29 22
rect 37 19 39 22
rect 55 19 57 22
rect -2 -40 0 13
rect 8 -40 10 13
rect 17 -10 19 13
rect 18 -14 19 -10
rect 17 -40 19 -14
rect 27 -40 29 13
rect 37 -40 39 13
rect 55 -40 57 13
rect -2 -47 0 -44
rect 8 -47 10 -44
rect 17 -47 19 -44
rect 27 -47 29 -44
rect 37 -47 39 -44
rect 55 -47 57 -44
<< polycontact >>
rect -6 0 -2 4
rect 4 -7 8 -3
rect 14 -14 18 -10
rect 23 -21 27 -17
rect 33 -28 37 -24
rect 51 -5 55 -1
<< metal1 >>
rect -13 31 73 35
rect -7 19 -3 31
rect 50 19 54 31
rect -17 0 -6 4
rect 41 -1 45 13
rect 58 -1 62 13
rect -17 -7 4 -3
rect 41 -5 51 -1
rect 58 -5 78 -1
rect -17 -14 14 -10
rect -17 -21 23 -17
rect -17 -28 33 -24
rect 41 -32 45 -5
rect 2 -36 45 -32
rect 2 -40 6 -36
rect 21 -40 25 -36
rect 41 -40 45 -36
rect 58 -40 62 -5
rect -7 -51 -3 -44
rect 11 -51 15 -44
rect 31 -51 35 -44
rect 50 -51 54 -44
rect -14 -55 73 -51
<< labels >>
rlabel metal1 -17 -7 8 -3 1 B
rlabel metal1 -17 0 -2 4 1 A
rlabel metal1 -17 -14 18 -10 1 C
rlabel metal1 -17 -21 27 -17 1 D
rlabel metal1 58 -5 78 -1 1 OUT
rlabel metal1 -13 31 73 35 5 VDD
rlabel metal1 41 -5 55 -1 1 5NOR
rlabel metal1 -14 -55 73 -51 1 GND
rlabel metal1 -17 -28 37 -24 1 E
<< end >>
