.include TSMC_180nm.txt

.param Supply=1.8
.param LAMBDA=0.09u
.param width_N=10*LAMBDA
.param width_P=20*LAMBDA
.global vdd gnd

Vdd vdd gnd 'SUPPLY'

vC cin gnd 0

vclk clk gnd pulse 0 1.8 0ns 0ns 0ns 5ns 10ns

vA0 a0 gnd pulse 0 1.8 0ns 0ns 0ns 10ns 20ns
vA1 a1 gnd pulse 0 1.8 0ns 0ns 0ns 15ns 30ns
vA2 a2 gnd pulse 0 1.8 0ns 0ns 0ns 20ns 40ns
vA3 a3 gnd pulse 0 1.8 0ns 0ns 0ns 25ns 50ns

vB0 b0 gnd pulse 0 1.8 0ns 0ns 0ns 10ns 20ns
vB1 b1 gnd pulse 0 1.8 0ns 0ns 0ns 15ns 30ns
vB2 b2 gnd pulse 0 1.8 0ns 0ns 0ns 20ns 40ns
vB3 b3 gnd pulse 0 1.8 0ns 0ns 0ns 25ns 50ns



* SPICE3 file created from nilavra_cla.ext - technology: scmos

.option scale=0.09u

M1000 3and_0/a_13_5# m1_n38_n151# m1_80_n107# 3and_0/w_0_n1# CMOSP w=6 l=2
+  ad=84 pd=52 as=108 ps=72
M1001 3and_0/a_13_n28# m1_n15_n136# m1_81_n168# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=40 ps=36
M1002 m1_89_n136# 3and_0/a_13_5# m1_81_n168# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 m1_80_n107# m1_n27_n143# 3and_0/a_13_5# 3and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 m1_89_n136# 3and_0/a_13_5# m1_80_n107# 3and_0/w_53_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1005 3and_0/a_13_5# m1_n15_n136# m1_80_n107# 3and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 3and_0/a_13_5# m1_n38_n151# 3and_0/a_23_n28# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1007 3and_0/a_23_n28# m1_n27_n143# 3and_0/a_13_n28# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 4or_0/a_0_n37# m1_156_n262# m1_191_n296# Gnd CMOSN w=4 l=2
+  ad=64 pd=48 as=92 ps=78
M1009 4or_0/a_0_n37# m1_178_n248# m1_191_n296# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 m1_271_n254# 4or_0/a_0_n37# m1_191_n296# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 4or_0/a_19_13# m1_156_n262# 4or_0/a_10_13# 4or_0/w_n13_7# CMOSP w=6 l=2
+  ad=48 pd=28 as=42 ps=26
M1012 m1_191_n296# m1_169_n255# 4or_0/a_0_n37# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 m1_271_n254# 4or_0/a_0_n37# m1_190_n221# 4or_0/w_n13_7# CMOSP w=6 l=2
+  ad=30 pd=22 as=60 ps=44
M1014 4or_0/a_0_13# m1_178_n248# m1_190_n221# 4or_0/w_n13_7# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1015 4or_0/a_0_n37# g2 4or_0/a_19_13# 4or_0/w_n13_7# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1016 4or_0/a_10_13# m1_169_n255# 4or_0/a_0_13# 4or_0/w_n13_7# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 m1_191_n296# g2 4or_0/a_0_n37# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 3and_1/a_13_5# m1_119_n93# m1_193_n48# 3and_1/w_0_n1# CMOSP w=6 l=2
+  ad=84 pd=52 as=108 ps=72
M1019 3and_1/a_13_n28# m1_n49_n10# m1_194_n109# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=40 ps=36
M1020 m1_276_n77# 3and_1/a_13_5# m1_194_n109# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1021 m1_193_n48# m1_n38_n95# 3and_1/a_13_5# 3and_1/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 m1_276_n77# 3and_1/a_13_5# m1_193_n48# 3and_1/w_53_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1023 3and_1/a_13_5# m1_n49_n10# m1_193_n48# 3and_1/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 3and_1/a_13_5# m1_119_n93# 3and_1/a_23_n28# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1025 3and_1/a_23_n28# m1_n38_n95# 3and_1/a_13_n28# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 3and_2/a_13_5# m1_322_n153# m1_393_n109# 3and_2/w_0_n1# CMOSP w=6 l=2
+  ad=84 pd=52 as=108 ps=72
M1027 3and_2/a_13_n28# g1 m1_467_n170# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=40 ps=36
M1028 m1_474_n138# 3and_2/a_13_5# m1_467_n170# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1029 m1_393_n109# m1_304_n147# 3and_2/a_13_5# 3and_2/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 m1_474_n138# 3and_2/a_13_5# m1_393_n109# 3and_2/w_53_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1031 3and_2/a_13_5# g1 m1_393_n109# 3and_2/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 3and_2/a_13_5# m1_322_n153# 3and_2/a_23_n28# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1033 3and_2/a_23_n28# m1_304_n147# 3and_2/a_13_n28# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 m1_65_79# p0 2and_0/a_13_5# 2and_0/w_0_n1# CMOSP w=6 l=2
+  ad=96 pd=68 as=48 ps=28
M1035 m1_69_49# 2and_0/a_13_5# 2and_0/a_6_n25# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1036 2and_0/a_13_5# c_in m1_65_79# 2and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 m1_69_49# 2and_0/a_13_5# m1_65_79# 2and_0/w_43_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1038 2and_0/a_13_5# p0 2and_0/a_13_n25# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1039 2and_0/a_13_n25# c_in 2and_0/a_6_n25# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 m1_71_n193# m1_n49_n231# 2and_1/a_13_5# 2and_1/w_0_n1# CMOSP w=6 l=2
+  ad=96 pd=68 as=48 ps=28
M1041 m1_79_n222# 2and_1/a_13_5# m1_72_n251# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1042 2and_1/a_13_5# m1_n38_n223# m1_71_n193# 2and_1/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 m1_79_n222# 2and_1/a_13_5# m1_71_n193# 2and_1/w_43_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1044 2and_1/a_13_5# m1_n49_n231# 2and_1/a_13_n25# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1045 2and_1/a_13_n25# m1_n38_n223# m1_72_n251# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 m1_192_n139# m1_119_n177# 2and_2/a_13_5# 2and_2/w_0_n1# CMOSP w=6 l=2
+  ad=96 pd=68 as=48 ps=28
M1047 2and_2/a_56_n25# 2and_2/a_13_5# m1_260_n199# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1048 2and_2/a_13_5# g1 m1_192_n139# 2and_2/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1049 2and_2/a_56_n25# 2and_2/a_13_5# m1_192_n139# 2and_2/w_43_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1050 2and_2/a_13_5# m1_119_n177# 2and_2/a_13_n25# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1051 2and_2/a_13_n25# g1 m1_260_n199# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 m1_391_n196# m1_322_n235# 2and_3/a_13_5# 2and_3/w_0_n1# CMOSP w=6 l=2
+  ad=96 pd=68 as=48 ps=28
M1053 m1_464_n225# 2and_3/a_13_5# m1_454_n254# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1054 2and_3/a_13_5# g2 m1_391_n196# 2and_3/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 m1_464_n225# 2and_3/a_13_5# m1_391_n196# 2and_3/w_43_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1056 2and_3/a_13_5# m1_322_n235# 2and_3/a_13_n25# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1057 2and_3/a_13_n25# g2 m1_454_n254# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 m1_478_n322# 5or_0/a_0_n44# m1_390_n290# 5or_0/w_n13_7# CMOSP w=6 l=2
+  ad=30 pd=22 as=60 ps=44
M1059 m1_471_n372# m1_347_n338# 5or_0/a_0_n44# Gnd CMOSN w=4 l=2
+  ad=100 pd=82 as=88 ps=68
M1060 m1_478_n322# 5or_0/a_0_n44# m1_471_n372# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1061 5or_0/a_0_n44# m1_357_n331# m1_471_n372# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 5or_0/a_0_n44# m1_376_n317# m1_471_n372# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 5or_0/a_19_13# m1_357_n331# 5or_0/a_10_13# 5or_0/w_n13_7# CMOSP w=6 l=2
+  ad=48 pd=28 as=42 ps=26
M1064 5or_0/a_0_13# m1_376_n317# m1_390_n290# 5or_0/w_n13_7# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1065 5or_0/a_29_13# m1_347_n338# 5or_0/a_19_13# 5or_0/w_n13_7# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1066 m1_471_n372# m1_366_n324# 5or_0/a_0_n44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 5or_0/a_10_13# m1_366_n324# 5or_0/a_0_13# 5or_0/w_n13_7# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 5or_0/a_0_n44# g3 5or_0/a_29_13# 5or_0/w_n13_7# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1069 5or_0/a_0_n44# g3 m1_471_n372# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 m1_60_n56# 2or_0/a_0_n30# m1_55_n22# 2or_0/w_n13_0# CMOSP w=6 l=2
+  ad=30 pd=22 as=60 ps=44
M1071 m1_57_n85# m1_4_n58# 2or_0/a_0_n30# Gnd CMOSN w=4 l=2
+  ad=60 pd=54 as=32 ps=24
M1072 2or_0/a_0_n30# m1_4_n58# 2or_0/a_0_6# 2or_0/w_n13_0# CMOSP w=6 l=2
+  ad=30 pd=22 as=48 ps=28
M1073 m1_60_n56# 2or_0/a_0_n30# m1_57_n85# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1074 2or_0/a_0_6# m1_n15_n51# m1_55_n22# 2or_0/w_n13_0# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 2or_0/a_0_n30# m1_n15_n51# m1_57_n85# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 m1_492_69# 5and_0/a_13_5# m1_394_98# 5and_0/w_73_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=156 ps=100
M1077 5and_0/a_13_5# m1_n38_n95# m1_394_98# 5and_0/w_0_n1# CMOSP w=6 l=2
+  ad=132 pd=80 as=0 ps=0
M1078 5and_0/a_43_n43# m1_304_46# 5and_0/a_33_n43# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1079 5and_0/a_33_n43# m1_n38_n95# 5and_0/a_23_n43# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1080 m1_394_98# m1_106_104# 5and_0/a_13_5# 5and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 5and_0/a_23_n43# m1_106_104# 5and_0/a_13_n43# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1082 m1_492_69# 5and_0/a_13_5# m1_488_22# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1083 5and_0/a_13_n43# c_in m1_488_22# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 5and_0/a_13_5# m1_322_39# m1_394_98# 5and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 5and_0/a_13_5# c_in m1_394_98# 5and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 m1_394_98# m1_304_46# 5and_0/a_13_5# 5and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 5and_0/a_13_5# m1_322_39# 5and_0/a_43_n43# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1088 m1_76_n307# 3or_0/a_0_n30# m1_71_n273# 3or_0/w_n13_7# CMOSP w=6 l=2
+  ad=30 pd=22 as=60 ps=44
M1089 m1_69_n343# m1_n11_n309# 3or_0/a_0_n30# Gnd CMOSN w=4 l=2
+  ad=68 pd=58 as=56 ps=44
M1090 m1_76_n307# 3or_0/a_0_n30# m1_69_n343# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1091 3or_0/a_0_n30# g1 3or_0/a_10_13# 3or_0/w_n13_7# CMOSP w=6 l=2
+  ad=36 pd=24 as=42 ps=26
M1092 3or_0/a_0_13# m1_n1_n302# m1_71_n273# 3or_0/w_n13_7# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1093 3or_0/a_10_13# m1_n11_n309# 3or_0/a_0_13# 3or_0/w_n13_7# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 3or_0/a_0_n30# g1 m1_69_n343# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 3or_0/a_0_n30# m1_n1_n302# m1_69_n343# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 4and_0/a_33_n36# m1_107_12# 4and_0/a_23_n36# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1097 4and_0/a_13_5# m1_107_12# m1_193_57# 4and_0/w_0_n1# CMOSP w=6 l=2
+  ad=96 pd=56 as=144 ps=96
M1098 4and_0/a_23_n36# m1_107_21# 4and_0/a_13_n36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1099 4and_0/a_13_n36# c_in m1_194_n12# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1100 m1_193_57# m1_107_21# 4and_0/a_13_5# 4and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 4and_0/a_13_5# c_in m1_193_57# 4and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 m1_271_28# 4and_0/a_13_5# m1_193_57# 4and_0/w_61_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 m1_271_28# 4and_0/a_13_5# m1_194_n12# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1104 m1_193_57# m1_119_6# 4and_0/a_13_5# 4and_0/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 4and_0/a_13_5# m1_119_6# 4and_0/a_33_n36# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1106 4and_1/a_33_n36# m1_304_n51# 4and_1/a_23_n36# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1107 4and_1/a_13_5# m1_304_n51# m1_393_n8# 4and_1/w_0_n1# CMOSP w=6 l=2
+  ad=96 pd=56 as=144 ps=96
M1108 4and_1/a_23_n36# m1_n38_n95# 4and_1/a_13_n36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1109 4and_1/a_13_n36# m1_346_n37# m1_476_n77# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1110 m1_393_n8# m1_n38_n95# 4and_1/a_13_5# 4and_1/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 4and_1/a_13_5# m1_346_n37# m1_393_n8# 4and_1/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 m1_483_n37# 4and_1/a_13_5# m1_393_n8# 4and_1/w_61_n1# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1113 m1_483_n37# 4and_1/a_13_5# m1_476_n77# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1114 m1_393_n8# m1_322_n59# 4and_1/a_13_5# 4and_1/w_0_n1# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 4and_1/a_13_5# m1_322_n59# 4and_1/a_33_n36# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
C0 5and_0/w_0_n1# m1_394_98# 0.08fF
C1 g1 m1_304_n147# 1.50fF
C2 m1_89_n136# m1_81_n168# 0.06fF
C3 m1_n1_n302# m2_n1_n302# 0.06fF
C4 m1_106_104# m5_55_n22# 0.07fF
C5 p1 m2_n38_n223# 0.08fF
C6 g1 m2_357_n331# 0.06fF
C7 m1_65_79# c_in 0.13fF
C8 m1_393_n8# m1_483_n37# 0.06fF
C9 g1 m1_n1_n302# 0.08fF
C10 m1_391_n196# m1_464_n225# 0.06fF
C11 2and_3/a_13_5# m1_454_n254# 0.02fF
C12 m1_n38_n95# m2_156_n262# 0.17fF
C13 5and_0/w_0_n1# c_in 0.08fF
C14 m1_357_n331# m1_347_n338# 1.01fF
C15 5or_0/w_n13_7# m1_390_n290# 0.06fF
C16 m1_366_n324# g3 0.08fF
C17 m1_n15_n136# m1_n27_n143# 0.57fF
C18 3and_0/w_0_n1# 3and_0/a_13_5# 0.05fF
C19 m1_60_n56# m5_55_n22# 0.05fF
C20 m2_107_n87# m4_57_n85# 0.15fF
C21 3and_1/a_13_5# m1_n38_n95# 0.16fF
C22 3or_0/w_n13_7# m1_n1_n302# 0.06fF
C23 m1_119_n93# m5_55_n22# 0.04fF
C24 4and_1/w_61_n1# m1_483_n37# 0.03fF
C25 m1_n38_n95# m2_n27_n143# 0.07fF
C26 m2_n15_n49# m2_n15_n136# 0.02fF
C27 m1_60_n56# m1_57_n85# 0.06fF
C28 m1_178_n248# m2_178_n248# 0.06fF
C29 4and_0/a_13_5# m1_194_n12# 0.02fF
C30 2and_2/w_0_n1# 2and_2/a_13_5# 0.02fF
C31 p0 m2_n27_n143# 0.12fF
C32 m1_190_n221# m5_55_n22# 0.01fF
C33 2or_0/a_0_n30# m1_55_n22# 0.04fF
C34 g1 g2 0.48fF
C35 carry2 m3_271_n254# 0.04fF
C36 m1_478_n322# m3_483_n421# 0.04fF
C37 m1_346_n37# m5_55_n22# 0.03fF
C38 m1_n49_n10# m2_n15_n49# 0.10fF
C39 m1_107_12# m1_119_6# 1.57fF
C40 4and_0/w_61_n1# m1_271_28# 0.03fF
C41 m1_107_21# 4and_0/a_13_5# 0.16fF
C42 g2 m2_119_n378# 0.16fF
C43 g2 m3_271_n254# 0.01fF
C44 p2 m2_119_n378# 0.15fF
C45 p2 m3_271_n254# 0.02fF
C46 g3 m4_57_n85# 0.05fF
C47 4and_0/w_0_n1# m1_107_21# 0.08fF
C48 m1_71_n193# m1_79_n222# 0.06fF
C49 2and_1/a_13_5# m1_72_n251# 0.02fF
C50 g0 m3_n69_48# 0.04fF
C51 m1_478_n322# m1_471_n372# 0.06fF
C52 g1 2and_2/w_0_n1# 0.08fF
C53 m1_474_n138# m2_366_n324# 0.06fF
C54 m1_322_n59# 4and_1/a_13_5# 0.12fF
C55 m1_454_n254# m5_55_n22# 0.02fF
C56 2and_1/w_0_n1# m1_71_n193# 0.06fF
C57 2and_1/w_43_n1# 2and_1/a_13_5# 0.08fF
C58 m1_107_12# m5_55_n22# 0.04fF
C59 3and_2/a_13_5# m1_393_n109# 0.13fF
C60 m1_71_n193# m5_55_n22# 0.03fF
C61 m1_72_n251# m4_57_n85# 0.03fF
C62 5or_0/a_0_n44# m1_471_n372# 0.33fF
C63 m1_390_n290# m1_478_n322# 0.06fF
C64 m1_178_n248# m1_156_n262# 0.08fF
C65 m2_376_n317# m5_55_n22# 0.07fF
C66 m1_178_n248# g2 0.08fF
C67 m1_71_n273# m1_76_n307# 0.06fF
C68 3or_0/a_0_n30# m1_69_n343# 0.21fF
C69 m1_n38_n95# m2_169_n255# 0.09fF
C70 5and_0/w_73_n1# 5and_0/a_13_5# 0.08fF
C71 m1_106_104# m1_304_46# 0.08fF
C72 c_in m1_322_39# 0.08fF
C73 3and_2/w_0_n1# 3and_2/a_13_5# 0.05fF
C74 5or_0/a_0_n44# m1_390_n290# 0.05fF
C75 m1_n11_n309# m2_n11_n309# 0.07fF
C76 m2_n11_n309# m4_57_n85# 0.16fF
C77 m1_n38_n95# m5_55_n22# 0.17fF
C78 4and_1/a_13_5# m1_476_n77# 0.02fF
C79 m2_156_n262# m2_169_n255# 0.18fF
C80 m1_57_n85# m1_n38_n95# 0.50fF
C81 m1_n15_n136# m1_n38_n151# 0.08fF
C82 3and_0/w_0_n1# m1_80_n107# 0.05fF
C83 3and_0/w_53_n1# 3and_0/a_13_5# 0.08fF
C84 m2_156_n262# m5_55_n22# 0.06fF
C85 5and_0/a_13_5# m1_488_22# 0.02fF
C86 m1_304_n147# m2_347_n338# 0.06fF
C87 g1 m2_304_n147# 0.09fF
C88 2and_2/a_13_5# 2and_2/a_56_n25# 0.05fF
C89 2and_0/w_43_n1# m1_69_49# 0.03fF
C90 p0 2and_0/a_13_5# 0.17fF
C91 g1 m3_145_n56# 0.09fF
C92 2and_0/w_0_n1# c_in 0.08fF
C93 m2_347_n338# m2_357_n331# 0.46fF
C94 m1_60_n56# m2_107_n87# 0.11fF
C95 m2_n49_n231# m2_n38_n223# 0.37fF
C96 m1_106_104# m2_n49_n231# 0.10fF
C97 5or_0/w_n13_7# m1_366_n324# 0.06fF
C98 m2_n15_n49# m4_57_n85# 0.09fF
C99 m2_n27_n143# m5_55_n22# 0.06fF
C100 m1_n49_n10# m2_119_n378# 0.07fF
C101 m1_193_57# m1_271_28# 0.06fF
C102 3and_1/a_13_5# m1_193_n48# 0.13fF
C103 2or_0/w_n13_0# m1_4_n58# 0.06fF
C104 m1_304_n51# m2_322_n393# 0.07fF
C105 m1_n15_n136# m2_n15_n136# 0.08fF
C106 g2 m2_347_n338# 0.06fF
C107 4or_0/a_0_n37# m1_271_n254# 0.05fF
C108 m1_346_n37# m2_n49_n231# 0.07fF
C109 g3 m3_94_n434# 0.01fF
C110 m1_119_6# m5_55_n22# 0.04fF
C111 m1_n38_n223# 2and_1/a_13_5# 0.04fF
C112 m1_169_n255# m1_156_n262# 0.86fF
C113 4or_0/w_n13_7# 4or_0/a_0_n37# 0.09fF
C114 m1_107_12# m2_107_n87# 0.06fF
C115 m1_169_n255# g2 0.08fF
C116 4and_1/w_0_n1# 4and_1/a_13_5# 0.05fF
C117 m1_346_n37# m1_304_n51# 0.08fF
C118 2and_3/w_0_n1# m1_322_n235# 0.08fF
C119 m1_393_n109# m5_55_n22# 0.05fF
C120 m1_n38_n95# m1_304_46# 1.45fF
C121 5and_0/w_73_n1# m1_394_98# 0.03fF
C122 g1 m1_322_n153# 0.08fF
C123 3and_2/w_0_n1# m1_393_n109# 0.05fF
C124 m2_169_n255# m5_55_n22# 0.06fF
C125 m2_n1_n302# m4_57_n85# 0.08fF
C126 m1_304_n147# m2_357_n331# 0.06fF
C127 3or_0/w_n13_7# m1_76_n307# 0.03fF
C128 m1_69_49# 2and_0/a_6_n25# 0.06fF
C129 g1 m4_57_n85# 0.17fF
C130 g1 m1_n11_n309# 0.77fF
C131 m1_n38_n95# m2_107_n87# 0.11fF
C132 5and_0/w_0_n1# m1_106_104# 0.08fF
C133 m1_357_n331# g3 0.08fF
C134 m1_366_n324# 5or_0/a_0_n44# 0.08fF
C135 m1_n27_n143# m1_n38_n151# 0.87fF
C136 m1_n15_n136# 3and_0/a_13_5# 0.04fF
C137 3and_0/w_53_n1# m1_80_n107# 0.03fF
C138 m2_119_n378# m4_57_n85# 0.42fF
C139 m1_119_n177# m1_260_n199# 0.03fF
C140 m3_271_n254# m4_57_n85# 0.10fF
C141 m3_178_n49# m5_55_n22# 0.14fF
C142 3or_0/w_n13_7# m1_n11_n309# 0.06fF
C143 m1_193_n48# m5_55_n22# 0.05fF
C144 m1_n38_n95# m2_n49_n231# 0.09fF
C145 c_in m3_n69_48# 0.08fF
C146 m2_n15_n136# m3_n69_48# 0.01fF
C147 2and_2/w_0_n1# m1_192_n139# 0.06fF
C148 2and_2/w_43_n1# 2and_2/a_13_5# 0.08fF
C149 m1_193_n48# m3_178_n49# 0.07fF
C150 p0 m2_n49_n231# 0.07fF
C151 m1_191_n296# m4_57_n85# 0.01fF
C152 m2_n27_n143# m2_107_n87# 0.03fF
C153 m1_n38_n95# m1_304_n51# 1.31fF
C154 c_in g0 0.04fF
C155 m1_89_n136# m2_n11_n309# 0.02fF
C156 m1_107_12# 4and_0/a_13_5# 0.08fF
C157 g2 m2_357_n331# 0.06fF
C158 m1_n49_n10# m3_n69_48# 0.01fF
C159 m2_n27_n143# m2_n49_n231# 0.22fF
C160 m1_n15_n51# m1_4_n58# 0.31fF
C161 3and_1/w_0_n1# m1_n49_n10# 0.08fF
C162 p3 m3_271_n254# 0.01fF
C163 carry0 m3_145_n56# 0.03fF
C164 carry1 m3_94_n434# 0.03fF
C165 4and_0/w_0_n1# m1_107_12# 0.08fF
C166 m1_190_n221# m1_271_n254# 0.06fF
C167 4or_0/a_0_n37# m1_191_n296# 0.25fF
C168 2and_3/a_13_5# m1_391_n196# 0.09fF
C169 2and_1/w_43_n1# m1_71_n193# 0.03fF
C170 m1_119_n177# m2_156_n262# 0.07fF
C171 5and_0/a_13_5# m1_394_98# 0.21fF
C172 m1_322_n153# m1_467_n170# 0.05fF
C173 3and_2/a_13_5# m1_474_n138# 0.05fF
C174 4or_0/w_n13_7# m1_190_n221# 0.06fF
C175 m1_156_n262# g2 1.02fF
C176 4and_1/w_0_n1# m1_393_n8# 0.08fF
C177 m1_n38_n223# m2_n38_n223# 0.08fF
C178 c_in 5and_0/a_13_5# 0.04fF
C179 m1_106_104# m1_322_39# 0.08fF
C180 3and_2/w_53_n1# 3and_2/a_13_5# 0.08fF
C181 m1_304_46# m5_55_n22# 0.02fF
C182 m1_322_39# m2_322_n393# 0.06fF
C183 5and_0/w_0_n1# m1_n38_n95# 0.08fF
C184 m1_347_n338# g3 1.27fF
C185 3and_0/w_53_n1# m1_89_n136# 0.03fF
C186 m1_n27_n143# 3and_0/a_13_5# 0.16fF
C187 m2_169_n255# m3_192_n139# 0.01fF
C188 m1_304_n147# m2_304_n147# 0.09fF
C189 g1 m2_322_n393# 0.07fF
C190 m1_322_n153# m2_347_n338# 0.06fF
C191 m1_192_n139# 2and_2/a_56_n25# 0.06fF
C192 2and_2/a_13_5# m1_260_n199# 0.02fF
C193 m3_192_n139# m5_55_n22# 0.05fF
C194 g1 m3_94_n434# 0.07fF
C195 m1_194_n109# m4_57_n85# 0.03fF
C196 2and_3/w_43_n1# m1_464_n225# 0.03fF
C197 m1_60_n56# m2_119_n378# 0.13fF
C198 5or_0/w_n13_7# m1_357_n331# 0.06fF
C199 m1_376_n317# m1_366_n324# 0.47fF
C200 m2_n49_n231# m5_55_n22# 0.06fF
C201 p1 m2_n49_n231# 0.09fF
C202 m1_119_n93# m2_119_n378# 0.09fF
C203 m1_65_79# m2_n27_n143# 0.07fF
C204 m1_391_n196# m5_55_n22# 0.02fF
C205 2or_0/a_0_n30# m1_60_n56# 0.05fF
C206 3and_1/a_13_5# m1_276_n77# 0.05fF
C207 m1_304_n51# m5_55_n22# 0.03fF
C208 m1_n49_n10# m1_55_n22# 0.44fF
C209 m1_119_6# 4and_0/a_13_5# 0.12fF
C210 m1_n15_n51# m2_n15_n49# 0.11fF
C211 m2_n27_n143# m2_n15_n49# 0.10fF
C212 2or_0/w_n13_0# 2or_0/a_0_n30# 0.09fF
C213 m1_322_n59# m2_322_n393# 0.08fF
C214 4and_0/w_0_n1# m1_119_6# 0.08fF
C215 m1_79_n222# m1_72_n251# 0.06fF
C216 m1_119_n177# m2_169_n255# 0.06fF
C217 m1_322_n235# m2_347_n338# 0.06fF
C218 g2 m2_304_n147# 0.07fF
C219 g2 m3_145_n56# 0.02fF
C220 m1_119_n177# m5_55_n22# 0.04fF
C221 p2 m2_304_n147# 0.05fF
C222 4and_1/a_13_5# m1_393_n8# 0.17fF
C223 p2 m3_145_n56# 0.02fF
C224 2and_1/w_43_n1# m1_79_n222# 0.03fF
C225 m1_n49_n231# 2and_1/a_13_5# 0.17fF
C226 m1_393_n109# m1_474_n138# 0.06fF
C227 m1_476_n77# m4_454_n254# 0.03fF
C228 m1_169_n255# 4or_0/a_0_n37# 0.08fF
C229 m1_346_n37# m1_322_n59# 0.08fF
C230 4and_1/w_61_n1# 4and_1/a_13_5# 0.08fF
C231 2and_3/w_0_n1# 2and_3/a_13_5# 0.02fF
C232 m1_467_n170# m4_454_n254# 0.03fF
C233 m2_357_n331# m2_366_n324# 0.35fF
C234 m1_n38_n95# m1_322_39# 0.17fF
C235 5and_0/w_73_n1# m1_492_69# 0.03fF
C236 m1_304_n147# m1_322_n153# 1.38fF
C237 g1 3and_2/a_13_5# 0.04fF
C238 3and_2/w_53_n1# m1_393_n109# 0.03fF
C239 m1_322_n153# m2_357_n331# 0.06fF
C240 m1_71_n273# m5_55_n22# 0.03fF
C241 3or_0/a_0_n30# m1_71_n273# 0.04fF
C242 m1_n38_n95# m2_119_n378# 0.19fF
C243 m1_492_69# m2_347_n338# 0.06fF
C244 c_in m2_n15_n136# 0.12fF
C245 m1_65_79# m5_55_n22# 0.03fF
C246 m1_357_n331# 5or_0/a_0_n44# 0.08fF
C247 m1_n38_n151# 3and_0/a_13_5# 0.12fF
C248 m1_492_69# m1_488_22# 0.06fF
C249 m1_276_n77# m2_169_n255# 0.06fF
C250 g1 m2_156_n262# 0.07fF
C251 m1_n1_n302# m1_n11_n309# 0.36fF
C252 2and_0/a_13_5# m1_65_79# 0.09fF
C253 m1_304_46# m2_n49_n231# 0.08fF
C254 5or_0/w_n13_7# m1_347_n338# 0.06fF
C255 m2_347_n338# m4_454_n254# 0.07fF
C256 m1_n49_n10# c_in 0.16fF
C257 m1_271_28# m1_194_n12# 0.06fF
C258 2and_2/w_43_n1# m1_192_n139# 0.03fF
C259 g2 m2_366_n324# 0.06fF
C260 2and_0/w_0_n1# p0 0.08fF
C261 m1_193_n48# m1_276_n77# 0.06fF
C262 m1_119_n93# m1_194_n109# 0.05fF
C263 m1_n38_n95# m1_322_n59# 0.17fF
C264 carry3 m3_483_n421# 0.04fF
C265 m1_471_n372# m4_57_n85# 0.01fF
C266 m1_322_n235# m2_357_n331# 0.06fF
C267 m1_n49_n10# m3_145_n56# 0.01fF
C268 g2 m4_57_n85# 0.09fF
C269 2and_3/w_0_n1# m5_55_n22# 0.06fF
C270 3and_1/w_0_n1# m1_119_n93# 0.08fF
C271 p2 m4_57_n85# 0.43fF
C272 m1_346_n37# m2_347_n338# 0.07fF
C273 m1_79_n222# m2_n1_n302# 0.07fF
C274 5and_0/a_13_5# m1_492_69# 0.05fF
C275 3and_2/a_13_5# m1_467_n170# 0.02fF
C276 m1_156_n262# 4or_0/a_0_n37# 0.08fF
C277 m1_119_6# m2_119_n378# 0.07fF
C278 c_in m1_107_21# 1.24fF
C279 4or_0/a_0_n37# g2 0.38fF
C280 4and_1/w_61_n1# m1_393_n8# 0.03fF
C281 g2 m1_322_n235# 0.78fF
C282 2and_1/w_0_n1# m1_n38_n223# 0.08fF
C283 m1_106_104# 5and_0/a_13_5# 0.16fF
C284 m1_322_39# m5_55_n22# 0.03fF
C285 g1 m2_169_n255# 0.06fF
C286 4and_1/w_0_n1# m1_346_n37# 0.08fF
C287 g1 m5_55_n22# 0.07fF
C288 g1 3or_0/a_0_n30# 0.30fF
C289 3and_2/w_0_n1# g1 0.08fF
C290 5and_0/w_0_n1# m1_304_46# 0.08fF
C291 2and_0/a_6_n25# m4_57_n85# 0.03fF
C292 m1_347_n338# 5or_0/a_0_n44# 0.08fF
C293 m2_357_n331# m4_454_n254# 0.07fF
C294 m1_304_n147# m2_322_n393# 0.07fF
C295 m3_483_n421# m4_454_n254# 0.11fF
C296 3or_0/w_n13_7# 3or_0/a_0_n30# 0.09fF
C297 m1_n38_n95# m2_347_n338# 0.07fF
C298 m1_376_n317# m1_357_n331# 0.08fF
C299 m2_304_n147# m4_57_n85# 0.07fF
C300 3and_1/w_0_n1# m1_n38_n95# 0.08fF
C301 m3_145_n56# m4_57_n85# 0.48fF
C302 2and_0/w_0_n1# 2and_0/a_13_5# 0.02fF
C303 m1_65_79# m2_n49_n231# 0.08fF
C304 m1_n49_n10# m4_57_n85# 0.09fF
C305 3and_1/a_13_5# m1_194_n109# 0.02fF
C306 m1_55_n22# m1_60_n56# 0.06fF
C307 2or_0/a_0_n30# m1_57_n85# 0.13fF
C308 m1_471_n372# m4_454_n254# 0.03fF
C309 m1_322_n59# m5_55_n22# 0.03fF
C310 m1_260_n199# m2_178_n248# 0.07fF
C311 3and_1/w_0_n1# 3and_1/a_13_5# 0.05fF
C312 m1_376_n317# m2_376_n317# 0.06fF
C313 m1_366_n324# m2_366_n324# 0.06fF
C314 2or_0/w_n13_0# m1_55_n22# 0.06fF
C315 m1_n38_n95# 4and_1/w_0_n1# 0.08fF
C316 m1_n15_n51# m3_n69_48# 0.01fF
C317 m2_n27_n143# m3_n69_48# 0.12fF
C318 p0 g0 0.19fF
C319 m1_n38_n151# m2_n38_n223# 0.09fF
C320 4and_0/w_0_n1# 4and_0/a_13_5# 0.05fF
C321 g2 m2_322_n393# 0.07fF
C322 m1_357_n331# m2_357_n331# 0.06fF
C323 g2 m3_94_n434# 0.01fF
C324 p3 m3_145_n56# 0.01fF
C325 p2 m3_94_n434# 0.02fF
C326 m1_194_n12# m4_57_n85# 0.03fF
C327 m1_193_57# m5_55_n22# 0.05fF
C328 m1_394_98# m1_492_69# 0.06fF
C329 m1_347_n338# m2_347_n338# 0.06fF
C330 m1_346_n37# 4and_1/a_13_5# 0.04fF
C331 2and_3/w_0_n1# m1_391_n196# 0.06fF
C332 2and_3/w_43_n1# 2and_3/a_13_5# 0.08fF
C333 m1_n27_n143# m2_n27_n143# 0.06fF
C334 3and_2/w_53_n1# m1_474_n138# 0.03fF
C335 m1_304_n147# 3and_2/a_13_5# 0.16fF
C336 m1_304_46# m1_322_39# 1.45fF
C337 m1_n38_n95# 5and_0/a_13_5# 0.08fF
C338 m1_76_n307# m4_57_n85# 0.04fF
C339 c_in m1_106_104# 0.68fF
C340 3and_0/a_13_5# m1_80_n107# 0.13fF
C341 2and_0/a_13_5# m1_69_49# 0.05fF
C342 m2_107_n87# m2_119_n378# 0.16fF
C343 m1_322_39# m2_n49_n231# 0.07fF
C344 5or_0/w_n13_7# g3 0.06fF
C345 m1_376_n317# m1_347_n338# 0.08fF
C346 m2_347_n338# m5_55_n22# 0.06fF
C347 2and_2/w_43_n1# 2and_2/a_56_n25# 0.03fF
C348 m1_119_n177# 2and_2/a_13_5# 0.17fF
C349 m1_322_n235# m2_366_n324# 0.06fF
C350 m1_n38_n95# 4and_1/a_13_5# 0.16fF
C351 m1_60_n56# m3_145_n56# 0.09fF
C352 m1_n49_n10# m1_60_n56# 0.17fF
C353 m1_169_n255# m2_169_n255# 0.06fF
C354 m1_119_n93# m3_145_n56# 0.01fF
C355 m1_4_n58# 2or_0/a_0_n30# 0.19fF
C356 m1_n49_n10# m1_119_n93# 0.08fF
C357 3and_1/w_0_n1# m1_193_n48# 0.05fF
C358 3and_1/w_53_n1# 3and_1/a_13_5# 0.08fF
C359 m1_156_n262# m2_156_n262# 0.06fF
C360 4and_0/w_61_n1# 4and_0/a_13_5# 0.08fF
C361 m1_192_n139# m5_55_n22# 0.05fF
C362 g1 m1_119_n177# 0.84fF
C363 g3 m3_271_n254# 0.01fF
C364 m1_119_n177# m2_119_n378# 0.10fF
C365 4or_0/w_n13_7# m1_271_n254# 0.03fF
C366 m1_271_28# m2_156_n262# 0.06fF
C367 c_in m1_107_12# 0.08fF
C368 m1_304_n51# m1_322_n59# 1.53fF
C369 g2 2and_3/a_13_5# 0.04fF
C370 2and_1/w_0_n1# m1_n49_n231# 0.08fF
C371 m1_n38_n223# m2_n11_n309# 0.07fF
C372 m2_n11_n309# m2_n1_n302# 0.11fF
C373 m2_169_n255# m2_178_n248# 0.11fF
C374 m2_366_n324# m4_454_n254# 0.08fF
C375 m2_178_n248# m5_55_n22# 0.09fF
C376 g1 m2_n11_n309# 0.02fF
C377 m1_304_n147# m5_55_n22# 0.02fF
C378 m1_n38_n95# m2_n15_n136# 0.08fF
C379 c_in m1_n38_n95# 0.08fF
C380 5and_0/w_0_n1# m1_322_39# 0.08fF
C381 3and_2/w_0_n1# m1_304_n147# 0.08fF
C382 g3 5or_0/a_0_n44# 0.48fF
C383 m1_n38_n151# m1_81_n168# 0.05fF
C384 3and_0/a_13_5# m1_89_n136# 0.05fF
C385 m2_357_n331# m5_55_n22# 0.05fF
C386 m1_322_n153# m2_322_n393# 0.08fF
C387 2and_2/a_56_n25# m1_260_n199# 0.06fF
C388 m1_76_n307# m3_94_n434# 0.02fF
C389 3or_0/w_n13_7# m1_71_n273# 0.06fF
C390 p0 2and_0/a_6_n25# 0.03fF
C391 p0 c_in 0.66fF
C392 m1_n38_n95# m2_304_n147# 0.11fF
C393 m1_366_n324# m1_357_n331# 0.92fF
C394 3and_0/w_0_n1# m1_n15_n136# 0.08fF
C395 m1_n38_n95# m3_145_n56# 0.09fF
C396 m1_60_n56# m4_57_n85# 0.06fF
C397 m2_322_n393# m4_57_n85# 0.07fF
C398 m1_55_n22# m5_55_n22# 0.03fF
C399 m1_n49_n10# m1_n38_n95# 1.46fF
C400 m3_94_n434# m4_57_n85# 0.12fF
C401 2and_0/w_0_n1# m1_65_79# 0.06fF
C402 2and_0/w_43_n1# 2and_0/a_13_5# 0.08fF
C403 m1_119_n93# m4_57_n85# 0.05fF
C404 m1_n15_n51# c_in 0.10fF
C405 c_in m2_n27_n143# 0.15fF
C406 m2_n27_n143# m2_n15_n136# 0.13fF
C407 m2_156_n262# m3_145_n56# 0.01fF
C408 m1_n49_n10# m2_156_n262# 0.07fF
C409 4and_0/a_13_5# m1_193_57# 0.17fF
C410 m1_271_n254# m3_271_n254# 0.02fF
C411 m2_n49_n231# m2_347_n338# 0.11fF
C412 g2 m5_55_n22# 0.04fF
C413 m1_n49_n10# 3and_1/a_13_5# 0.04fF
C414 3and_1/w_53_n1# m1_193_n48# 0.03fF
C415 m1_483_n37# m1_476_n77# 0.06fF
C416 m1_464_n225# m1_454_n254# 0.06fF
C417 m2_n49_n231# m3_n69_48# 0.13fF
C418 m1_390_n290# m5_55_n22# 0.02fF
C419 m1_4_n58# m3_n69_48# 0.04fF
C420 m1_n49_n10# m2_n27_n143# 0.09fF
C421 m1_107_21# m1_107_12# 1.60fF
C422 4and_0/w_0_n1# m1_193_57# 0.08fF
C423 m1_322_n235# m2_322_n393# 0.08fF
C424 p3 m2_322_n393# 0.08fF
C425 m1_464_n225# m2_376_n317# 0.06fF
C426 m1_260_n199# m4_57_n85# 0.03fF
C427 m1_271_n254# m1_191_n296# 0.06fF
C428 m1_304_n51# m2_347_n338# 0.07fF
C429 g1 2and_2/a_13_5# 0.04fF
C430 p3 m3_94_n434# 0.01fF
C431 g0 m2_n49_n231# 0.09fF
C432 2and_1/a_13_5# m1_71_n193# 0.09fF
C433 m2_366_n324# m2_376_n317# 0.10fF
C434 m1_474_n138# m1_467_n170# 0.06fF
C435 m1_192_n139# m3_192_n139# 0.04fF
C436 4or_0/a_0_n37# m1_190_n221# 0.04fF
C437 c_in m1_119_6# 0.08fF
C438 2and_3/w_43_n1# m1_391_n196# 0.03fF
C439 m1_76_n307# m1_69_n343# 0.06fF
C440 m1_304_46# 5and_0/a_13_5# 0.08fF
C441 m1_322_n153# 3and_2/a_13_5# 0.12fF
C442 4or_0/w_n13_7# m1_178_n248# 0.06fF
C443 m1_394_98# m5_55_n22# 0.05fF
C444 4and_1/w_0_n1# m1_304_n51# 0.08fF
C445 m1_69_n343# m4_57_n85# 0.03fF
C446 5or_0/w_n13_7# m1_478_n322# 0.03fF
C447 3and_0/a_13_5# m1_81_n168# 0.02fF
C448 m1_80_n107# m1_89_n136# 0.06fF
C449 m1_107_21# m2_n27_n143# 0.11fF
C450 m1_n38_n95# m4_57_n85# 0.11fF
C451 c_in m5_55_n22# 0.15fF
C452 g1 m2_119_n378# 0.13fF
C453 m1_65_79# m1_69_49# 0.06fF
C454 2and_0/a_13_5# 2and_0/a_6_n25# 0.02fF
C455 g1 3or_0/w_n13_7# 0.06fF
C456 m1_n49_n231# m2_n49_n231# 0.07fF
C457 g1 m3_271_n254# 0.07fF
C458 m1_322_n235# m1_454_n254# 0.03fF
C459 2and_3/a_13_5# m1_464_n225# 0.05fF
C460 2and_0/a_13_5# c_in 0.04fF
C461 m1_376_n317# g3 0.08fF
C462 m1_366_n324# m1_347_n338# 0.08fF
C463 5or_0/w_n13_7# 5or_0/a_0_n44# 0.09fF
C464 3and_0/w_0_n1# m1_n27_n143# 0.08fF
C465 m2_156_n262# m4_57_n85# 0.15fF
C466 m1_n49_n10# m5_55_n22# 0.11fF
C467 m1_69_49# m2_n15_n49# 0.09fF
C468 m1_276_n77# m1_194_n109# 0.06fF
C469 m1_393_n8# m5_55_n22# 0.05fF
C470 m1_119_6# m1_194_n12# 0.04fF
C471 2or_0/w_n13_0# m1_60_n56# 0.03fF
C472 m2_n15_n49# m3_n69_48# 0.13fF
C473 m1_80_n107# m1_n38_n95# 0.82fF
C474 m1_107_21# m1_119_6# 0.08fF
C475 4and_0/w_61_n1# m1_193_57# 0.03fF
C476 m1_81_n168# m4_57_n85# 0.04fF
C477 m1_n49_n231# m1_72_n251# 0.03fF
C478 2and_1/a_13_5# m1_79_n222# 0.05fF
C479 m1_304_n51# 4and_1/a_13_5# 0.08fF
C480 m1_322_n235# 2and_3/a_13_5# 0.17fF
C481 m1_454_n254# m4_454_n254# 0.03fF
C482 m1_107_21# m5_55_n22# 0.04fF
C483 m1_483_n37# m2_357_n331# 0.06fF
C484 2and_1/w_0_n1# 2and_1/a_13_5# 0.02fF
C485 m1_n49_n231# m2_n11_n309# 0.07fF
C486 m1_79_n222# m4_57_n85# 0.04fF
C487 5or_0/a_0_n44# m1_478_n322# 0.05fF
C488 4or_0/w_n13_7# m1_169_n255# 0.06fF
C489 m2_376_n317# m4_454_n254# 0.07fF
C490 m2_366_n324# m5_55_n22# 0.05fF
C491 3or_0/a_0_n30# m1_76_n307# 0.05fF
C492 m1_322_n153# m5_55_n22# 0.03fF
C493 m1_n38_n95# m2_n38_n223# 0.10fF
C494 5and_0/w_0_n1# 5and_0/a_13_5# 0.08fF
C495 m1_106_104# m1_n38_n95# 0.81fF
C496 c_in m1_304_46# 0.08fF
C497 3and_2/w_0_n1# m1_322_n153# 0.08fF
C498 m2_169_n255# m4_57_n85# 0.07fF
C499 m4_57_n85# m5_55_n22# 1.21fF
C500 m1_n11_n309# 3or_0/a_0_n30# 0.08fF
C501 4and_1/a_13_5# m1_483_n37# 0.05fF
C502 m1_322_n59# m1_476_n77# 0.04fF
C503 m1_n38_n95# m2_322_n393# 0.12fF
C504 m1_304_46# m2_304_n147# 0.08fF
C505 3and_0/w_0_n1# m1_n38_n151# 0.08fF
C506 m1_57_n85# m4_57_n85# 0.03fF
C507 m1_322_39# m1_488_22# 0.05fF
C508 g1 m2_347_n338# 0.06fF
C509 2and_2/a_13_5# m1_192_n139# 0.09fF
C510 m1_119_n93# m1_n38_n95# 1.47fF
C511 2and_0/w_43_n1# m1_65_79# 0.03fF
C512 c_in m2_n49_n231# 0.34fF
C513 m2_n27_n143# m2_n38_n223# 0.18fF
C514 m1_106_104# m2_n27_n143# 0.11fF
C515 m1_4_n58# c_in 0.02fF
C516 5or_0/w_n13_7# m1_376_n317# 0.06fF
C517 m1_119_n93# m2_156_n262# 0.07fF
C518 m1_n49_n10# m2_107_n87# 0.07fF
C519 4and_0/a_13_5# m1_271_28# 0.05fF
C520 2and_2/w_0_n1# m1_119_n177# 0.08fF
C521 m1_322_n235# m5_55_n22# 0.04fF
C522 m1_119_n93# 3and_1/a_13_5# 0.12fF
C523 3and_1/w_53_n1# m1_276_n77# 0.03fF
C524 m1_n38_n95# m1_346_n37# 0.92fF
C525 m1_n49_n10# m2_n49_n231# 0.12fF
C526 m1_80_n107# m5_55_n22# 0.03fF
C527 2or_0/w_n13_0# m1_n15_n51# 0.06fF
C528 m1_322_n59# m2_347_n338# 0.07fF
C529 m1_304_n51# m2_304_n147# 0.09fF
C530 m1_271_n254# g2 0.03fF
C531 c_in 4and_0/a_13_5# 0.04fF
C532 g3 m3_145_n56# 0.01fF
C533 m1_n38_n223# m1_n49_n231# 0.68fF
C534 m1_322_39# 5and_0/a_13_5# 0.12fF
C535 m1_119_n177# m3_145_n56# 0.01fF
C536 4or_0/w_n13_7# m1_156_n262# 0.06fF
C537 m1_178_n248# m1_169_n255# 0.44fF
C538 c_in 4and_0/w_0_n1# 0.08fF
C539 4or_0/w_n13_7# g2 0.06fF
C540 4and_1/w_0_n1# m1_322_n59# 0.08fF
C541 2and_3/w_0_n1# g2 0.08fF
C542 m5_55_n22# Gnd 0.28fF **FLOATING
C543 m4_57_n85# Gnd 0.23fF **FLOATING
C544 m3_483_n421# Gnd 0.07fF **FLOATING
C545 m3_192_n139# Gnd 0.00fF **FLOATING
C546 m3_94_n434# Gnd 0.12fF **FLOATING
C547 m2_376_n317# Gnd 0.42fF **FLOATING
C548 m2_366_n324# Gnd 0.48fF **FLOATING
C549 m2_n11_n309# Gnd 0.11fF **FLOATING
C550 m2_n38_n223# Gnd 0.64fF **FLOATING
C551 m2_n15_n136# Gnd 0.30fF **FLOATING
C552 m2_357_n331# Gnd 0.57fF **FLOATING
C553 m2_119_n378# Gnd 0.81fF **FLOATING
C554 m2_107_n87# Gnd 0.11fF **FLOATING
C555 m2_156_n262# Gnd 0.11fF **FLOATING
C556 m2_322_n393# Gnd 0.91fF **FLOATING
C557 m2_304_n147# Gnd 0.25fF **FLOATING
C558 m2_347_n338# Gnd 0.71fF **FLOATING
C559 m2_n49_n231# Gnd 1.42fF **FLOATING
C560 m2_n27_n143# Gnd 0.19fF **FLOATING
C561 carry3 Gnd 0.09fF **FLOATING
C562 carry2 Gnd 0.06fF **FLOATING
C563 carry0 Gnd 0.05fF **FLOATING
C564 carry1 Gnd 0.05fF **FLOATING
C565 p3 Gnd 0.38fF **FLOATING
C566 p2 Gnd 0.41fF **FLOATING
C567 p1 Gnd 0.29fF **FLOATING
C568 g0 Gnd 0.05fF **FLOATING
C569 m1_476_n77# Gnd 0.39fF
C570 m1_483_n37# Gnd 0.14fF
C571 m1_393_n8# Gnd 0.38fF
C572 4and_1/a_13_5# Gnd 0.52fF
C573 m1_322_n59# Gnd 0.29fF
C574 m1_304_n51# Gnd 0.40fF
C575 m1_346_n37# Gnd 0.48fF
C576 4and_1/w_61_n1# Gnd 0.43fF
C577 4and_1/w_0_n1# Gnd 0.99fF
C578 m1_194_n12# Gnd 0.34fF
C579 m1_271_28# Gnd 0.23fF
C580 m1_193_57# Gnd 0.25fF
C581 4and_0/a_13_5# Gnd 0.52fF
C582 m1_119_6# Gnd 0.64fF
C583 m1_107_12# Gnd 0.65fF
C584 m1_107_21# Gnd 0.62fF
C585 4and_0/w_61_n1# Gnd 0.43fF
C586 4and_0/w_0_n1# Gnd 0.99fF
C587 m1_69_n343# Gnd 0.13fF
C588 m1_76_n307# Gnd 0.26fF
C589 m1_71_n273# Gnd 0.31fF
C590 3or_0/a_0_n30# Gnd 0.46fF
C591 m1_n11_n309# Gnd 0.34fF
C592 m1_n1_n302# Gnd 0.29fF
C593 3or_0/w_n13_7# Gnd 1.21fF
C594 m1_488_22# Gnd 0.41fF
C595 m1_492_69# Gnd 0.14fF
C596 m1_394_98# Gnd 0.42fF
C597 5and_0/a_13_5# Gnd 0.62fF
C598 m1_322_39# Gnd 0.69fF
C599 m1_304_46# Gnd 0.37fF
C600 m1_n38_n95# Gnd 1.16fF
C601 m1_106_104# Gnd 1.75fF
C602 5and_0/w_73_n1# Gnd 0.43fF
C603 5and_0/w_0_n1# Gnd 1.18fF
C604 m1_57_n85# Gnd 0.31fF
C605 m1_55_n22# Gnd 0.28fF
C606 2or_0/a_0_n30# Gnd 0.35fF
C607 m1_4_n58# Gnd 0.29fF
C608 m1_n15_n51# Gnd 0.23fF
C609 2or_0/w_n13_0# Gnd 1.03fF
C610 m1_471_n372# Gnd 0.42fF
C611 m1_478_n322# Gnd 0.25fF
C612 m1_390_n290# Gnd 0.31fF
C613 5or_0/a_0_n44# Gnd 0.65fF
C614 g3 Gnd 0.86fF
C615 m1_347_n338# Gnd 0.61fF
C616 m1_357_n331# Gnd 0.55fF
C617 m1_366_n324# Gnd 0.51fF
C618 m1_376_n317# Gnd 0.45fF
C619 5or_0/w_n13_7# Gnd 1.55fF
C620 m1_454_n254# Gnd 0.33fF
C621 m1_464_n225# Gnd 0.17fF
C622 m1_391_n196# Gnd 0.28fF
C623 2and_3/a_13_5# Gnd 0.37fF
C624 m1_322_n235# Gnd 0.53fF
C625 g2 Gnd 1.04fF
C626 2and_3/w_43_n1# Gnd 0.43fF
C627 2and_3/w_0_n1# Gnd 0.67fF
C628 m1_260_n199# Gnd 0.31fF
C629 2and_2/a_56_n25# Gnd 0.11fF
C630 m1_192_n139# Gnd 0.28fF
C631 2and_2/a_13_5# Gnd 0.37fF
C632 m1_119_n177# Gnd 0.52fF
C633 2and_2/w_43_n1# Gnd 0.43fF
C634 2and_2/w_0_n1# Gnd 0.67fF
C635 m1_72_n251# Gnd 0.33fF
C636 m1_79_n222# Gnd 0.17fF
C637 m1_71_n193# Gnd 0.36fF
C638 2and_1/a_13_5# Gnd 0.37fF
C639 m1_n49_n231# Gnd 0.51fF
C640 m1_n38_n223# Gnd 0.46fF
C641 2and_1/w_43_n1# Gnd 0.43fF
C642 2and_1/w_0_n1# Gnd 0.67fF
C643 2and_0/a_6_n25# Gnd 0.29fF
C644 m1_69_49# Gnd 0.17fF
C645 m1_65_79# Gnd 0.69fF
C646 2and_0/a_13_5# Gnd 0.37fF
C647 p0 Gnd 0.17fF
C648 2and_0/w_43_n1# Gnd 0.43fF
C649 2and_0/w_0_n1# Gnd 0.67fF
C650 m1_467_n170# Gnd 0.37fF
C651 m1_474_n138# Gnd 0.17fF
C652 m1_393_n109# Gnd 0.33fF
C653 3and_2/a_13_5# Gnd 0.43fF
C654 m1_322_n153# Gnd 0.46fF
C655 m1_304_n147# Gnd 0.59fF
C656 g1 Gnd 1.40fF
C657 3and_2/w_53_n1# Gnd 0.43fF
C658 3and_2/w_0_n1# Gnd 0.83fF
C659 m1_194_n109# Gnd 0.32fF
C660 m1_276_n77# Gnd 0.18fF
C661 m1_193_n48# Gnd 0.06fF
C662 3and_1/a_13_5# Gnd 0.43fF
C663 m1_119_n93# Gnd 0.57fF
C664 m1_n49_n10# Gnd 0.45fF
C665 3and_1/w_53_n1# Gnd 0.43fF
C666 3and_1/w_0_n1# Gnd 0.83fF
C667 m1_191_n296# Gnd 0.36fF
C668 m1_271_n254# Gnd 0.23fF
C669 m1_190_n221# Gnd 0.28fF
C670 4or_0/a_0_n37# Gnd 0.54fF
C671 m1_156_n262# Gnd 0.51fF
C672 m1_169_n255# Gnd 0.37fF
C673 m1_178_n248# Gnd 0.31fF
C674 4or_0/w_n13_7# Gnd 1.39fF
C675 m1_81_n168# Gnd 0.36fF
C676 m1_89_n136# Gnd 0.14fF
C677 m1_80_n107# Gnd 0.39fF
C678 3and_0/a_13_5# Gnd 0.43fF
C679 m1_n38_n151# Gnd 0.43fF
C680 m1_n27_n143# Gnd 0.37fF
C681 m1_n15_n136# Gnd 0.29fF
C682 3and_0/w_53_n1# Gnd 0.43fF
C683 3and_0/w_0_n1# Gnd 0.83fF
