magic
tech scmos
timestamp 1638764848
<< metal1 >>
rect 106 104 369 111
rect -100 81 15 86
rect 65 79 73 87
rect 364 66 369 104
rect 394 98 402 106
rect 382 69 400 74
rect 492 69 503 73
rect 498 68 503 69
rect 193 57 201 65
rect 364 62 399 66
rect 340 55 392 59
rect -108 49 -42 53
rect -31 50 8 53
rect -38 49 8 50
rect 69 49 90 53
rect -69 48 -63 49
rect -49 47 -42 49
rect 81 48 90 49
rect 304 47 407 52
rect 304 46 311 47
rect -60 40 -1 44
rect 322 40 403 44
rect 322 39 328 40
rect 129 28 202 32
rect 271 28 293 32
rect 288 27 293 28
rect 107 21 195 25
rect 488 22 496 29
rect 107 14 199 18
rect 107 12 113 14
rect 119 7 196 11
rect 119 6 126 7
rect -49 -10 79 -3
rect 55 -22 63 -14
rect -15 -51 2 -47
rect -103 -58 -38 -54
rect -31 -58 -8 -54
rect 4 -58 14 -54
rect -102 -73 -31 -67
rect 73 -73 79 -10
rect 194 -12 201 -6
rect 393 -8 401 0
rect 346 -33 353 -30
rect 346 -37 403 -33
rect 483 -37 491 -33
rect 486 -38 491 -37
rect 193 -48 201 -40
rect 340 -44 396 -40
rect 304 -47 311 -44
rect 304 -51 403 -47
rect 322 -58 398 -54
rect 322 -59 328 -58
rect 73 -77 194 -73
rect 276 -77 292 -73
rect 476 -77 484 -70
rect 287 -78 292 -77
rect 57 -85 63 -78
rect 107 -84 193 -80
rect 107 -87 113 -84
rect -38 -90 -31 -88
rect 107 -90 112 -87
rect -38 -95 112 -90
rect 119 -91 197 -87
rect 119 -93 126 -91
rect 80 -107 88 -99
rect 106 -109 112 -95
rect 194 -109 201 -103
rect 393 -109 401 -101
rect -15 -136 5 -132
rect 89 -136 97 -132
rect -27 -139 -21 -137
rect 192 -139 200 -131
rect 299 -138 398 -134
rect 474 -138 486 -134
rect -27 -143 3 -139
rect 480 -140 486 -138
rect -38 -146 -31 -144
rect 304 -145 392 -141
rect -38 -150 4 -146
rect 304 -147 311 -145
rect -38 -151 -31 -150
rect 322 -152 398 -148
rect 322 -153 328 -152
rect 81 -168 87 -161
rect 136 -168 197 -164
rect 467 -170 475 -163
rect 119 -177 214 -173
rect 71 -193 79 -185
rect 193 -197 200 -191
rect 260 -199 268 -193
rect 391 -196 399 -188
rect -38 -218 -31 -216
rect -38 -223 15 -218
rect 79 -222 97 -218
rect 190 -221 198 -213
rect -49 -227 -42 -224
rect 284 -225 395 -221
rect 464 -225 480 -221
rect -49 -231 17 -227
rect 178 -244 183 -243
rect 72 -251 78 -244
rect 178 -248 191 -244
rect 169 -251 174 -250
rect 169 -255 196 -251
rect 271 -254 278 -249
rect 156 -258 162 -256
rect 156 -262 197 -258
rect 71 -273 79 -265
rect 111 -269 197 -265
rect -1 -298 5 -296
rect -1 -302 9 -298
rect 94 -303 100 -302
rect -11 -309 5 -305
rect 76 -307 100 -303
rect -102 -313 7 -312
rect -102 -316 -11 -313
rect -5 -316 7 -313
rect 69 -343 75 -336
rect 111 -356 116 -269
rect 191 -296 198 -290
rect 284 -356 290 -225
rect 474 -227 480 -225
rect 322 -234 396 -230
rect 322 -235 328 -234
rect 454 -254 461 -248
rect 390 -290 398 -282
rect 376 -313 382 -311
rect 376 -317 391 -313
rect 366 -320 371 -319
rect 366 -324 393 -320
rect 478 -322 488 -318
rect 357 -327 362 -326
rect 357 -331 391 -327
rect 347 -334 352 -333
rect 347 -338 391 -334
rect -103 -362 290 -356
rect 346 -345 392 -341
rect -103 -378 311 -371
rect -103 -393 328 -387
rect 346 -401 353 -345
rect 391 -373 398 -367
rect 471 -372 478 -366
rect -103 -407 353 -401
rect 94 -448 100 -428
rect 146 -448 152 -430
rect 272 -451 279 -423
rect 483 -435 488 -413
<< m2contact >>
rect 376 69 382 74
rect 335 55 340 60
rect -38 50 -31 55
rect 123 28 129 33
rect -38 -58 -31 -51
rect 60 -56 66 -50
rect 335 -44 340 -39
rect 106 -117 112 -109
rect 294 -139 299 -134
rect 130 -169 136 -164
rect -11 -319 -5 -313
rect 130 -351 136 -344
<< metal2 >>
rect -38 129 382 136
rect -38 55 -31 129
rect -38 -51 -31 50
rect 123 33 129 129
rect 376 74 382 129
rect 335 -39 340 55
rect 66 -56 149 -50
rect 335 -112 340 -44
rect 112 -117 340 -112
rect -11 -346 -5 -319
rect 130 -344 136 -169
rect -11 -351 130 -346
rect 294 -346 299 -139
rect 136 -351 299 -346
<< m3contact >>
rect 106 104 114 111
rect -49 47 -42 53
rect -49 -10 -42 -3
rect 81 44 90 53
rect -27 39 -21 44
rect 498 68 503 73
rect 304 46 311 52
rect 322 39 328 44
rect 107 22 113 29
rect 288 27 293 32
rect 107 12 113 18
rect 119 6 126 11
rect 346 -37 353 -30
rect 486 -38 491 -33
rect -15 -49 -8 -43
rect -15 -62 -8 -55
rect 304 -51 311 -44
rect 322 -59 328 -54
rect -38 -73 -31 -67
rect 287 -78 292 -73
rect 107 -87 113 -80
rect -38 -95 -31 -88
rect 119 -93 126 -87
rect -15 -136 -8 -130
rect -27 -143 -21 -137
rect 91 -138 97 -132
rect -38 -151 -31 -144
rect 119 -179 126 -173
rect -38 -223 -31 -216
rect 91 -224 97 -218
rect -49 -231 -42 -224
rect -1 -302 5 -296
rect -11 -309 -5 -303
rect 260 -199 268 -193
rect 178 -248 183 -243
rect 169 -255 174 -250
rect 156 -262 162 -256
rect 480 -140 486 -134
rect 304 -147 311 -141
rect 322 -153 328 -148
rect 474 -227 480 -221
rect 322 -235 328 -230
rect 376 -317 382 -311
rect 366 -324 371 -319
rect 357 -331 362 -326
rect 347 -338 352 -333
rect 119 -378 126 -371
rect 322 -393 328 -387
<< metal3 >>
rect -49 118 353 123
rect -49 117 122 118
rect 306 117 353 118
rect -49 53 -42 117
rect -49 -3 -42 47
rect -49 -224 -42 -10
rect -27 105 106 111
rect -27 44 -21 105
rect -38 -88 -31 -73
rect -38 -144 -31 -95
rect -27 -137 -21 39
rect 81 16 90 44
rect 107 29 113 104
rect -15 9 90 16
rect -15 -43 -8 9
rect -15 -130 -8 -62
rect 107 -80 113 12
rect 119 -87 126 6
rect 288 -28 293 27
rect 156 -34 293 -28
rect -38 -216 -31 -151
rect 91 -174 97 -138
rect -11 -180 97 -174
rect 119 -173 126 -93
rect -11 -303 -5 -180
rect 91 -256 97 -224
rect -1 -262 97 -256
rect -1 -296 5 -262
rect 119 -371 126 -179
rect 156 -256 162 -34
rect 178 -49 199 -43
rect 304 -44 311 46
rect 287 -121 292 -78
rect 169 -126 292 -121
rect 169 -250 174 -126
rect 192 -139 197 -133
rect 304 -141 311 -51
rect 260 -200 268 -199
rect 178 -205 268 -200
rect 178 -243 183 -205
rect 304 -378 311 -147
rect 322 -54 328 39
rect 346 -30 353 117
rect 498 8 503 68
rect 357 2 503 8
rect 322 -148 328 -59
rect 357 -81 363 2
rect 322 -230 328 -153
rect 322 -387 328 -235
rect 347 -87 363 -81
rect 347 -333 352 -87
rect 486 -93 491 -38
rect 357 -98 491 -93
rect 357 -326 362 -98
rect 486 -99 491 -98
rect 480 -179 486 -140
rect 366 -184 486 -179
rect 366 -319 371 -184
rect 474 -267 480 -227
rect 376 -274 480 -267
rect 376 -311 382 -274
<< m4contact >>
rect -69 48 -63 53
rect -4 -59 1 -54
rect 145 -56 152 -50
rect 94 -307 100 -302
rect 271 -254 278 -249
rect 483 -322 488 -317
rect 483 -421 488 -414
rect 94 -434 100 -428
rect 146 -437 152 -430
rect 272 -432 279 -423
<< metal4 >>
rect -69 3 -63 48
rect -69 -2 1 3
rect -4 -54 1 -2
rect 94 -428 100 -307
rect 146 -430 152 -56
rect 272 -249 278 -248
rect 272 -423 278 -254
rect 483 -414 488 -322
<< m5contact >>
rect 66 20 72 27
rect 488 22 496 29
rect 194 -12 201 -6
rect 57 -85 63 -78
rect 81 -168 87 -161
rect 72 -251 78 -244
rect 69 -343 75 -336
rect 476 -77 484 -70
rect 194 -109 201 -103
rect 467 -170 475 -163
rect 193 -197 200 -191
rect 454 -254 461 -248
rect 191 -296 198 -290
rect 391 -373 398 -367
rect 471 -372 478 -366
<< metal5 >>
rect 66 5 72 20
rect 66 -1 89 5
rect 84 -7 89 -1
rect 84 -12 194 -7
rect 84 -64 89 -12
rect 488 -23 493 22
rect 488 -28 503 -23
rect 57 -70 143 -64
rect 57 -78 63 -70
rect 136 -104 143 -70
rect 498 -72 503 -28
rect 484 -77 503 -72
rect 136 -109 194 -104
rect 136 -148 143 -109
rect 83 -154 143 -148
rect 83 -161 89 -154
rect 87 -168 89 -161
rect 83 -204 89 -168
rect 498 -164 503 -77
rect 475 -170 503 -164
rect 143 -197 193 -192
rect 143 -204 147 -197
rect 83 -210 147 -204
rect 83 -246 89 -210
rect 78 -251 89 -246
rect 83 -338 89 -251
rect 498 -250 503 -170
rect 461 -254 503 -250
rect 457 -255 503 -254
rect 191 -338 197 -296
rect 75 -343 197 -338
rect 191 -368 197 -343
rect 191 -372 391 -368
rect 498 -367 503 -255
rect 478 -372 503 -367
<< m6contact >>
rect 394 98 402 106
rect 65 79 73 87
rect 193 57 201 65
rect 393 -8 401 0
rect 55 -22 63 -14
rect 193 -48 201 -40
rect 80 -107 88 -99
rect 393 -109 401 -101
rect 192 -139 200 -131
rect 71 -193 79 -185
rect 391 -196 399 -188
rect 190 -221 198 -213
rect 71 -273 79 -265
rect 390 -290 398 -282
<< metal6 >>
rect 386 98 394 106
rect 386 87 392 98
rect 73 82 392 87
rect 94 -15 99 82
rect 63 -20 99 -15
rect 94 -99 99 -20
rect 88 -107 99 -99
rect 93 -122 99 -107
rect 178 64 183 82
rect 178 57 193 64
rect 178 -40 184 57
rect 387 0 392 82
rect 387 -8 393 0
rect 178 -48 193 -40
rect 178 -49 201 -48
rect 93 -127 106 -122
rect 101 -185 106 -127
rect 79 -190 106 -185
rect 101 -265 106 -190
rect 178 -131 184 -49
rect 387 -101 392 -8
rect 387 -109 393 -101
rect 178 -139 192 -131
rect 178 -213 184 -139
rect 387 -188 392 -109
rect 387 -196 391 -188
rect 178 -221 190 -213
rect 79 -271 106 -265
rect 387 -282 393 -196
rect 387 -290 390 -282
use 2and  2and_0
timestamp 1638596035
transform 1 0 4 0 1 56
box -5 -36 71 30
use 4and  4and_0
timestamp 1638596374
transform 1 0 195 0 1 35
box -5 -47 89 30
use 5and  5and_0
timestamp 1638596562
transform 1 0 395 0 1 76
box -5 -54 101 30
use 2or  2or_0
timestamp 1638596115
transform 1 0 16 0 1 -44
box -17 -41 49 28
use 3and  3and_0
timestamp 1638596191
transform 1 0 8 0 1 -129
box -5 -39 81 30
use 3and  3and_1
timestamp 1638596191
transform 1 0 195 0 1 -70
box -5 -39 81 30
use 4and  4and_1
timestamp 1638596374
transform 1 0 395 0 1 -30
box -5 -47 89 30
use 2and  2and_1
timestamp 1638596035
transform 1 0 8 0 1 -215
box -5 -36 71 30
use 2and  2and_2
timestamp 1638596035
transform 1 0 194 0 1 -161
box -5 -36 71 30
use 3and  3and_2
timestamp 1638596191
transform 1 0 395 0 1 -131
box -5 -39 81 30
use 3or  3or_0
timestamp 1638596283
transform 1 0 20 0 1 -302
box -17 -41 59 35
use 4or  4or_0
timestamp 1638596467
transform 1 0 205 0 1 -248
box -17 -48 69 35
use 2and  2and_3
timestamp 1638596035
transform 1 0 393 0 1 -218
box -5 -36 71 30
use 5or  5or_0
timestamp 1638596680
transform 1 0 405 0 1 -317
box -17 -55 78 35
<< labels >>
rlabel metal1 -60 40 -51 44 1 p0
rlabel metal1 94 -448 100 -437 1 carry1
rlabel metal1 146 -448 152 -439 1 carry0
rlabel metal1 272 -451 279 -440 1 carry2
rlabel metal1 483 -435 488 -424 1 carry3
rlabel metal1 -103 -407 -92 -401 1 g3
rlabel metal1 -103 -393 -92 -387 1 p3
rlabel metal1 -103 -378 -92 -371 1 p2
rlabel metal1 -103 -362 -92 -356 1 g2
rlabel metal1 -102 -316 -93 -312 1 g1
rlabel metal1 -102 -73 -87 -67 1 p1
rlabel metal1 -103 -58 -86 -54 1 c_in
rlabel metal1 -108 49 -89 53 1 g0
<< end >>
