* SPICE3 file created from dflipflop.ext - technology: scmos

.option scale=0.09u

M1000 a_403_429# a_358_341# a_320_399# w_390_423# pfet w=50 l=2
+  ad=250 pd=110 as=1250 ps=540
M1001 a_320_399# a_332_489# a_365_399# w_352_393# pfet w=80 l=2
+  ad=0 pd=0 as=480 ps=172
M1002 a_365_341# a_320_364# a_358_341# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=200 ps=90
M1003 a_327_364# a_324_489# a_320_364# Gnd nfet w=20 l=2
+  ad=600 pd=280 as=100 ps=50
M1004 a_403_429# a_332_489# a_403_374# Gnd nfet w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1005 a_327_364# a_332_489# a_365_341# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_403_374# a_358_341# a_327_364# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_433_403# a_403_429# a_320_399# w_420_431# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1008 a_327_399# a_324_489# a_320_399# w_314_393# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1009 a_320_364# a_332_489# a_327_399# w_314_393# pfet w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1010 a_365_399# a_320_364# a_358_341# w_352_393# pfet w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1011 a_433_403# a_403_429# a_327_364# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 a_320_399# a_327_399# 0.82fF
C1 a_320_399# w_420_431# 0.11fF
C2 a_403_374# a_403_429# 0.41fF
C3 a_327_399# a_320_364# 0.82fF
C4 a_358_341# w_352_393# 0.20fF
C5 a_332_489# w_314_393# 0.08fF
C6 a_358_341# a_332_489# 0.58fF
C7 a_320_399# a_324_489# 0.01fF
C8 a_320_399# a_365_399# 0.82fF
C9 a_332_489# w_352_393# 0.08fF
C10 a_327_364# a_403_374# 0.44fF
C11 a_433_403# w_420_431# 0.06fF
C12 a_324_489# a_320_364# 0.06fF
C13 a_403_429# a_332_489# 0.06fF
C14 a_358_341# a_327_364# 0.05fF
C15 a_320_399# w_314_393# 0.25fF
C16 a_358_341# a_320_399# 0.85fF
C17 a_358_341# w_390_423# 0.08fF
C18 a_320_399# w_352_393# 0.25fF
C19 a_320_364# w_314_393# 0.10fF
C20 a_327_364# a_403_429# 0.29fF
C21 a_320_399# a_332_489# 0.02fF
C22 a_358_341# a_320_364# 0.72fF
C23 a_320_399# a_403_429# 0.54fF
C24 a_332_489# w_390_423# 0.36fF
C25 a_320_364# w_352_393# 0.17fF
C26 a_332_489# a_320_364# 0.47fF
C27 a_403_429# w_390_423# 0.07fF
C28 a_358_341# a_365_341# 0.47fF
C29 a_403_429# a_433_403# 0.05fF
C30 a_327_399# w_314_393# 0.01fF
C31 a_327_364# a_320_364# 0.26fF
C32 a_320_399# w_390_423# 0.16fF
C33 a_327_364# a_433_403# 0.21fF
C34 a_320_399# a_320_364# 0.09fF
C35 a_324_489# w_314_393# 0.08fF
C36 a_320_399# a_433_403# 0.45fF
C37 a_358_341# a_365_399# 0.82fF
C38 a_327_364# a_365_341# 0.41fF
C39 a_403_429# w_420_431# 0.06fF
C40 a_324_489# a_332_489# 0.17fF
C41 a_365_399# w_352_393# 0.01fF
C42 a_403_374# Gnd 0.01fF
C43 a_365_341# Gnd 0.01fF
C44 a_327_364# Gnd 0.86fF
C45 a_433_403# Gnd 0.09fF
C46 a_403_429# Gnd 0.24fF
C47 a_320_399# Gnd 0.64fF
C48 a_358_341# Gnd 0.63fF
C49 a_320_364# Gnd 0.60fF
C50 a_332_489# Gnd 0.74fF
C51 a_324_489# Gnd 0.17fF
C52 w_420_431# Gnd 1.25fF
C53 w_390_423# Gnd 1.49fF
C54 w_352_393# Gnd 2.96fF
C55 w_314_393# Gnd 2.96fF
