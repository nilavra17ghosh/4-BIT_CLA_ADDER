magic
tech scmos
timestamp 1732021772
<< nwell >>
rect 314 393 346 485
rect 352 393 384 485
rect 390 423 414 485
rect 420 431 444 483
<< ntransistor >>
rect 325 364 327 384
rect 363 341 365 381
rect 371 341 373 381
rect 401 374 403 414
rect 409 374 411 414
rect 431 403 433 423
<< ptransistor >>
rect 325 399 327 479
rect 333 399 335 479
rect 363 399 365 479
rect 371 399 373 479
rect 401 429 403 479
rect 431 437 433 477
<< ndiffusion >>
rect 324 364 325 384
rect 327 364 328 384
rect 362 341 363 381
rect 365 341 366 381
rect 370 341 371 381
rect 373 341 374 381
rect 400 374 401 414
rect 403 374 404 414
rect 408 374 409 414
rect 411 374 412 414
rect 430 403 431 423
rect 433 403 434 423
<< pdiffusion >>
rect 324 399 325 479
rect 327 399 328 479
rect 332 399 333 479
rect 335 399 336 479
rect 362 399 363 479
rect 365 399 366 479
rect 370 399 371 479
rect 373 399 374 479
rect 400 429 401 479
rect 403 429 404 479
rect 430 437 431 477
rect 433 437 434 477
<< ndcontact >>
rect 320 364 324 384
rect 328 364 332 384
rect 358 341 362 381
rect 366 341 370 381
rect 374 341 378 381
rect 396 374 400 414
rect 404 374 408 414
rect 412 374 416 414
rect 426 403 430 423
rect 434 403 438 423
<< pdcontact >>
rect 320 399 324 479
rect 328 399 332 479
rect 336 399 340 479
rect 358 399 362 479
rect 366 399 370 479
rect 374 399 378 479
rect 396 429 400 479
rect 404 429 408 479
rect 426 437 430 477
rect 434 437 438 477
<< polysilicon >>
rect 325 479 327 489
rect 333 479 335 489
rect 363 479 365 489
rect 371 479 373 489
rect 401 479 403 489
rect 401 414 403 429
rect 409 414 411 489
rect 431 477 433 480
rect 431 423 433 437
rect 325 384 327 399
rect 333 392 335 399
rect 363 381 365 399
rect 371 381 373 399
rect 325 361 327 364
rect 431 400 433 403
rect 401 371 403 374
rect 409 371 411 374
rect 363 338 365 341
rect 371 338 373 341
<< polycontact >>
rect 324 489 328 493
rect 332 489 336 493
rect 362 489 366 493
rect 370 489 374 493
rect 400 489 404 493
rect 408 489 412 493
rect 427 426 431 430
<< metal1 >>
rect 332 500 412 504
rect 324 493 328 497
rect 332 493 336 500
rect 348 493 366 497
rect 323 480 324 486
rect 320 479 324 480
rect 336 390 340 399
rect 348 390 352 493
rect 370 493 374 500
rect 384 493 404 497
rect 374 480 376 484
rect 374 479 379 480
rect 320 387 352 390
rect 358 389 362 399
rect 384 389 388 493
rect 408 493 412 500
rect 396 481 400 484
rect 423 481 444 486
rect 391 480 400 481
rect 396 479 400 480
rect 426 477 430 481
rect 408 430 416 432
rect 408 429 427 430
rect 412 426 427 429
rect 434 429 438 437
rect 412 414 416 426
rect 434 425 449 429
rect 434 423 438 425
rect 320 384 324 387
rect 358 384 388 389
rect 328 332 332 364
rect 358 381 362 384
rect 374 339 378 341
rect 426 394 430 403
rect 420 390 444 394
rect 396 368 400 374
rect 420 368 423 390
rect 396 364 423 368
rect 396 339 400 364
rect 374 335 400 339
rect 374 332 378 335
rect 328 328 378 332
<< m2contact >>
rect 318 480 323 486
rect 376 480 381 485
rect 391 481 396 487
rect 417 481 423 487
<< metal2 >>
rect 323 485 391 486
rect 323 482 376 485
rect 381 482 391 485
rect 396 482 417 486
use project1_inverter  project1_inverter_0
timestamp 1731863481
transform 1 0 91 0 1 53
box 0 0 1 1
<< end >>
