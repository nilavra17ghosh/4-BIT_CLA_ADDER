magic
tech scmos
timestamp 1732107157
<< nwell >>
rect 1301 -732 1333 -640
rect 1339 -732 1371 -640
rect 1377 -702 1401 -640
rect 1407 -694 1431 -642
rect 1503 -695 1528 -672
rect 220 -752 310 -734
rect -315 -868 -283 -776
rect -277 -868 -245 -776
rect -239 -838 -215 -776
rect -209 -830 -185 -778
rect -120 -888 -88 -796
rect -82 -888 -50 -796
rect -44 -858 -20 -796
rect -14 -850 10 -798
rect 220 -844 310 -826
rect 908 -857 973 -839
rect 981 -857 1005 -839
rect 517 -877 554 -859
rect 560 -877 584 -859
rect 708 -898 763 -880
rect 769 -898 793 -880
rect 220 -936 310 -918
rect 1091 -920 1181 -902
rect 1304 -922 1336 -830
rect 1342 -922 1374 -830
rect 1380 -892 1404 -830
rect 1410 -884 1434 -832
rect 1503 -885 1528 -862
rect -317 -1059 -285 -967
rect -279 -1059 -247 -967
rect -241 -1029 -217 -967
rect -211 -1021 -187 -969
rect 516 -976 573 -958
rect 908 -963 963 -945
rect 969 -963 993 -945
rect -119 -1071 -87 -979
rect -81 -1071 -49 -979
rect -43 -1041 -19 -979
rect -13 -1033 11 -981
rect 708 -1003 754 -985
rect 761 -1003 785 -985
rect 220 -1029 310 -1011
rect 1091 -1018 1181 -1000
rect 521 -1062 567 -1044
rect 574 -1062 598 -1044
rect 908 -1064 954 -1046
rect 961 -1064 985 -1046
rect 707 -1094 744 -1076
rect 750 -1094 774 -1076
rect 230 -1133 267 -1115
rect 273 -1133 297 -1115
rect 1091 -1118 1181 -1100
rect 1302 -1111 1334 -1019
rect 1340 -1111 1372 -1019
rect 1378 -1081 1402 -1019
rect 1408 -1073 1432 -1021
rect 1502 -1074 1527 -1051
rect 521 -1148 558 -1130
rect 564 -1148 588 -1130
rect 906 -1151 943 -1133
rect 949 -1151 973 -1133
rect -317 -1253 -285 -1161
rect -279 -1253 -247 -1161
rect -241 -1223 -217 -1161
rect -211 -1215 -187 -1163
rect -115 -1253 -83 -1161
rect -77 -1253 -45 -1161
rect -39 -1223 -15 -1161
rect -9 -1215 15 -1163
rect 705 -1173 782 -1155
rect 229 -1208 266 -1190
rect 272 -1208 296 -1190
rect 520 -1227 587 -1209
rect 1091 -1216 1181 -1198
rect 905 -1242 991 -1224
rect 229 -1283 266 -1265
rect 272 -1283 296 -1265
rect 1303 -1300 1335 -1208
rect 1341 -1300 1373 -1208
rect 1379 -1270 1403 -1208
rect 1409 -1262 1433 -1210
rect 1500 -1263 1525 -1240
rect -317 -1437 -285 -1345
rect -279 -1437 -247 -1345
rect -241 -1407 -217 -1345
rect -211 -1399 -187 -1347
rect -112 -1435 -80 -1343
rect -74 -1435 -42 -1343
rect -36 -1405 -12 -1343
rect -6 -1397 18 -1345
rect 229 -1358 266 -1340
rect 272 -1358 296 -1340
rect 1304 -1488 1336 -1396
rect 1342 -1488 1374 -1396
rect 1380 -1458 1404 -1396
rect 1410 -1450 1434 -1398
rect 1503 -1451 1528 -1428
<< ntransistor >>
rect 1312 -761 1314 -741
rect 231 -792 233 -788
rect 247 -792 249 -788
rect 257 -792 259 -788
rect 267 -792 269 -788
rect 277 -792 279 -788
rect -304 -897 -302 -877
rect -266 -920 -264 -880
rect -258 -920 -256 -880
rect -228 -887 -226 -847
rect -220 -887 -218 -847
rect -198 -858 -196 -838
rect 1350 -784 1352 -744
rect 1358 -784 1360 -744
rect 1388 -751 1390 -711
rect 1396 -751 1398 -711
rect 1418 -722 1420 -702
rect 1515 -707 1517 -703
rect 297 -792 299 -788
rect -109 -917 -107 -897
rect -71 -940 -69 -900
rect -63 -940 -61 -900
rect -33 -907 -31 -867
rect -25 -907 -23 -867
rect -3 -878 -1 -858
rect 231 -884 233 -880
rect 247 -884 249 -880
rect 257 -884 259 -880
rect 267 -884 269 -880
rect 277 -884 279 -880
rect 297 -884 299 -880
rect 528 -901 530 -897
rect 538 -901 540 -897
rect 571 -901 573 -897
rect 919 -899 921 -895
rect 929 -899 931 -895
rect 939 -899 941 -895
rect 949 -899 951 -895
rect 959 -899 961 -895
rect 992 -899 994 -895
rect 719 -933 721 -929
rect 729 -933 731 -929
rect 739 -933 741 -929
rect 749 -933 751 -929
rect 780 -933 782 -929
rect -306 -1088 -304 -1068
rect -268 -1111 -266 -1071
rect -260 -1111 -258 -1071
rect -230 -1078 -228 -1038
rect -222 -1078 -220 -1038
rect -200 -1049 -198 -1029
rect 231 -976 233 -972
rect 247 -976 249 -972
rect 257 -976 259 -972
rect 267 -976 269 -972
rect 277 -976 279 -972
rect 297 -976 299 -972
rect 1102 -960 1104 -956
rect 1118 -960 1120 -956
rect 1128 -960 1130 -956
rect 1138 -960 1140 -956
rect 1148 -960 1150 -956
rect 1315 -951 1317 -931
rect 1168 -960 1170 -956
rect 1353 -974 1355 -934
rect 1361 -974 1363 -934
rect 1391 -941 1393 -901
rect 1399 -941 1401 -901
rect 1421 -912 1423 -892
rect 1515 -897 1517 -893
rect 527 -1006 529 -1002
rect 537 -1006 539 -1002
rect 555 -1006 557 -1002
rect -108 -1100 -106 -1080
rect -70 -1123 -68 -1083
rect -62 -1123 -60 -1083
rect -32 -1090 -30 -1050
rect -24 -1090 -22 -1050
rect -2 -1061 0 -1041
rect 919 -998 921 -994
rect 929 -998 931 -994
rect 939 -998 941 -994
rect 949 -998 951 -994
rect 980 -998 982 -994
rect 719 -1030 721 -1026
rect 729 -1030 731 -1026
rect 739 -1030 741 -1026
rect 772 -1030 774 -1026
rect 231 -1069 233 -1065
rect 247 -1069 249 -1065
rect 257 -1069 259 -1065
rect 267 -1069 269 -1065
rect 277 -1069 279 -1065
rect 297 -1069 299 -1065
rect 1102 -1058 1104 -1054
rect 1118 -1058 1120 -1054
rect 1128 -1058 1130 -1054
rect 1138 -1058 1140 -1054
rect 1148 -1058 1150 -1054
rect 532 -1089 534 -1085
rect 542 -1089 544 -1085
rect 552 -1089 554 -1085
rect 585 -1089 587 -1085
rect 1168 -1058 1170 -1054
rect 919 -1091 921 -1087
rect 929 -1091 931 -1087
rect 939 -1091 941 -1087
rect 972 -1091 974 -1087
rect 718 -1118 720 -1114
rect 728 -1118 730 -1114
rect 761 -1118 763 -1114
rect 241 -1157 243 -1153
rect 251 -1157 253 -1153
rect 284 -1157 286 -1153
rect -306 -1282 -304 -1262
rect -268 -1305 -266 -1265
rect -260 -1305 -258 -1265
rect -230 -1272 -228 -1232
rect -222 -1272 -220 -1232
rect -200 -1243 -198 -1223
rect 532 -1172 534 -1168
rect 542 -1172 544 -1168
rect 575 -1172 577 -1168
rect -104 -1282 -102 -1262
rect -66 -1305 -64 -1265
rect -58 -1305 -56 -1265
rect -28 -1272 -26 -1232
rect -20 -1272 -18 -1232
rect 2 -1243 4 -1223
rect 1313 -1140 1315 -1120
rect 1102 -1158 1104 -1154
rect 1118 -1158 1120 -1154
rect 1128 -1158 1130 -1154
rect 1138 -1158 1140 -1154
rect 1148 -1158 1150 -1154
rect 1168 -1158 1170 -1154
rect 1351 -1163 1353 -1123
rect 1359 -1163 1361 -1123
rect 1389 -1130 1391 -1090
rect 1397 -1130 1399 -1090
rect 1419 -1101 1421 -1081
rect 1514 -1086 1516 -1082
rect 917 -1175 919 -1171
rect 927 -1175 929 -1171
rect 960 -1175 962 -1171
rect 716 -1217 718 -1213
rect 726 -1217 728 -1213
rect 735 -1217 737 -1213
rect 745 -1217 747 -1213
rect 764 -1217 766 -1213
rect 240 -1232 242 -1228
rect 250 -1232 252 -1228
rect 283 -1232 285 -1228
rect 531 -1264 533 -1260
rect 541 -1264 543 -1260
rect 550 -1264 552 -1260
rect 569 -1264 571 -1260
rect 1102 -1256 1104 -1252
rect 1118 -1256 1120 -1252
rect 1128 -1256 1130 -1252
rect 1138 -1256 1140 -1252
rect 1148 -1256 1150 -1252
rect 1168 -1256 1170 -1252
rect 916 -1293 918 -1289
rect 926 -1293 928 -1289
rect 935 -1293 937 -1289
rect 945 -1293 947 -1289
rect 955 -1293 957 -1289
rect 973 -1293 975 -1289
rect 240 -1307 242 -1303
rect 250 -1307 252 -1303
rect 283 -1307 285 -1303
rect 1314 -1329 1316 -1309
rect -306 -1466 -304 -1446
rect -268 -1489 -266 -1449
rect -260 -1489 -258 -1449
rect -230 -1456 -228 -1416
rect -222 -1456 -220 -1416
rect -200 -1427 -198 -1407
rect 1352 -1352 1354 -1312
rect 1360 -1352 1362 -1312
rect 1390 -1319 1392 -1279
rect 1398 -1319 1400 -1279
rect 1420 -1290 1422 -1270
rect 1512 -1275 1514 -1271
rect 240 -1382 242 -1378
rect 250 -1382 252 -1378
rect 283 -1382 285 -1378
rect -101 -1464 -99 -1444
rect -63 -1487 -61 -1447
rect -55 -1487 -53 -1447
rect -25 -1454 -23 -1414
rect -17 -1454 -15 -1414
rect 5 -1425 7 -1405
rect 1315 -1517 1317 -1497
rect 1353 -1540 1355 -1500
rect 1361 -1540 1363 -1500
rect 1391 -1507 1393 -1467
rect 1399 -1507 1401 -1467
rect 1421 -1478 1423 -1458
rect 1515 -1463 1517 -1459
<< ptransistor >>
rect 1312 -726 1314 -646
rect 1320 -726 1322 -646
rect 1350 -726 1352 -646
rect 1358 -726 1360 -646
rect 1388 -696 1390 -646
rect 1418 -688 1420 -648
rect 1515 -688 1517 -680
rect 231 -746 233 -740
rect 247 -746 249 -740
rect 257 -746 259 -740
rect 267 -746 269 -740
rect 277 -746 279 -740
rect 297 -746 299 -740
rect -304 -862 -302 -782
rect -296 -862 -294 -782
rect -266 -862 -264 -782
rect -258 -862 -256 -782
rect -228 -832 -226 -782
rect -198 -824 -196 -784
rect -109 -882 -107 -802
rect -101 -882 -99 -802
rect -71 -882 -69 -802
rect -63 -882 -61 -802
rect -33 -852 -31 -802
rect -3 -844 -1 -804
rect 231 -838 233 -832
rect 247 -838 249 -832
rect 257 -838 259 -832
rect 267 -838 269 -832
rect 277 -838 279 -832
rect 297 -838 299 -832
rect 919 -851 921 -845
rect 929 -851 931 -845
rect 939 -851 941 -845
rect 949 -851 951 -845
rect 959 -851 961 -845
rect 992 -851 994 -845
rect 528 -871 530 -865
rect 538 -871 540 -865
rect 571 -871 573 -865
rect 719 -892 721 -886
rect 729 -892 731 -886
rect 739 -892 741 -886
rect 749 -892 751 -886
rect 780 -892 782 -886
rect 231 -930 233 -924
rect 247 -930 249 -924
rect 257 -930 259 -924
rect 267 -930 269 -924
rect 277 -930 279 -924
rect 297 -930 299 -924
rect -306 -1053 -304 -973
rect -298 -1053 -296 -973
rect -268 -1053 -266 -973
rect -260 -1053 -258 -973
rect -230 -1023 -228 -973
rect 1102 -914 1104 -908
rect 1118 -914 1120 -908
rect 1128 -914 1130 -908
rect 1138 -914 1140 -908
rect 1148 -914 1150 -908
rect 1168 -914 1170 -908
rect 919 -957 921 -951
rect 929 -957 931 -951
rect 939 -957 941 -951
rect 949 -957 951 -951
rect 980 -957 982 -951
rect 1315 -916 1317 -836
rect 1323 -916 1325 -836
rect 1353 -916 1355 -836
rect 1361 -916 1363 -836
rect 1391 -886 1393 -836
rect 1421 -878 1423 -838
rect 1515 -878 1517 -870
rect -200 -1015 -198 -975
rect -108 -1065 -106 -985
rect -100 -1065 -98 -985
rect -70 -1065 -68 -985
rect -62 -1065 -60 -985
rect -32 -1035 -30 -985
rect 527 -970 529 -964
rect 537 -970 539 -964
rect 555 -970 557 -964
rect -2 -1027 0 -987
rect 719 -997 721 -991
rect 729 -997 731 -991
rect 739 -997 741 -991
rect 772 -997 774 -991
rect 231 -1023 233 -1017
rect 247 -1023 249 -1017
rect 257 -1023 259 -1017
rect 267 -1023 269 -1017
rect 277 -1023 279 -1017
rect 297 -1023 299 -1017
rect 1102 -1012 1104 -1006
rect 1118 -1012 1120 -1006
rect 1128 -1012 1130 -1006
rect 1138 -1012 1140 -1006
rect 1148 -1012 1150 -1006
rect 1168 -1012 1170 -1006
rect 532 -1056 534 -1050
rect 542 -1056 544 -1050
rect 552 -1056 554 -1050
rect 585 -1056 587 -1050
rect 919 -1058 921 -1052
rect 929 -1058 931 -1052
rect 939 -1058 941 -1052
rect 972 -1058 974 -1052
rect 718 -1088 720 -1082
rect 728 -1088 730 -1082
rect 761 -1088 763 -1082
rect 1102 -1112 1104 -1106
rect 1118 -1112 1120 -1106
rect 1128 -1112 1130 -1106
rect 1138 -1112 1140 -1106
rect 1148 -1112 1150 -1106
rect 1168 -1112 1170 -1106
rect 241 -1127 243 -1121
rect 251 -1127 253 -1121
rect 284 -1127 286 -1121
rect 532 -1142 534 -1136
rect 542 -1142 544 -1136
rect 575 -1142 577 -1136
rect -306 -1247 -304 -1167
rect -298 -1247 -296 -1167
rect -268 -1247 -266 -1167
rect -260 -1247 -258 -1167
rect -230 -1217 -228 -1167
rect -200 -1209 -198 -1169
rect -104 -1247 -102 -1167
rect -96 -1247 -94 -1167
rect -66 -1247 -64 -1167
rect -58 -1247 -56 -1167
rect -28 -1217 -26 -1167
rect 917 -1145 919 -1139
rect 927 -1145 929 -1139
rect 960 -1145 962 -1139
rect 716 -1167 718 -1161
rect 726 -1167 728 -1161
rect 735 -1167 737 -1161
rect 745 -1167 747 -1161
rect 764 -1167 766 -1161
rect 2 -1209 4 -1169
rect 240 -1202 242 -1196
rect 250 -1202 252 -1196
rect 283 -1202 285 -1196
rect 1313 -1105 1315 -1025
rect 1321 -1105 1323 -1025
rect 1351 -1105 1353 -1025
rect 1359 -1105 1361 -1025
rect 1389 -1075 1391 -1025
rect 1419 -1067 1421 -1027
rect 1514 -1067 1516 -1059
rect 1102 -1210 1104 -1204
rect 1118 -1210 1120 -1204
rect 1128 -1210 1130 -1204
rect 1138 -1210 1140 -1204
rect 1148 -1210 1150 -1204
rect 1168 -1210 1170 -1204
rect 531 -1221 533 -1215
rect 541 -1221 543 -1215
rect 550 -1221 552 -1215
rect 569 -1221 571 -1215
rect 916 -1236 918 -1230
rect 926 -1236 928 -1230
rect 935 -1236 937 -1230
rect 945 -1236 947 -1230
rect 955 -1236 957 -1230
rect 973 -1236 975 -1230
rect 240 -1277 242 -1271
rect 250 -1277 252 -1271
rect 283 -1277 285 -1271
rect 1314 -1294 1316 -1214
rect 1322 -1294 1324 -1214
rect 1352 -1294 1354 -1214
rect 1360 -1294 1362 -1214
rect 1390 -1264 1392 -1214
rect 1420 -1256 1422 -1216
rect 1512 -1256 1514 -1248
rect -306 -1431 -304 -1351
rect -298 -1431 -296 -1351
rect -268 -1431 -266 -1351
rect -260 -1431 -258 -1351
rect -230 -1401 -228 -1351
rect -200 -1393 -198 -1353
rect -101 -1429 -99 -1349
rect -93 -1429 -91 -1349
rect -63 -1429 -61 -1349
rect -55 -1429 -53 -1349
rect -25 -1399 -23 -1349
rect 5 -1391 7 -1351
rect 240 -1352 242 -1346
rect 250 -1352 252 -1346
rect 283 -1352 285 -1346
rect 1315 -1482 1317 -1402
rect 1323 -1482 1325 -1402
rect 1353 -1482 1355 -1402
rect 1361 -1482 1363 -1402
rect 1391 -1452 1393 -1402
rect 1421 -1444 1423 -1404
rect 1515 -1444 1517 -1436
<< ndiffusion >>
rect 1311 -761 1312 -741
rect 1314 -761 1315 -741
rect 230 -792 231 -788
rect 233 -792 234 -788
rect 246 -792 247 -788
rect 249 -792 257 -788
rect 259 -792 261 -788
rect 265 -792 267 -788
rect 269 -792 277 -788
rect 279 -792 280 -788
rect -305 -897 -304 -877
rect -302 -897 -301 -877
rect -267 -920 -266 -880
rect -264 -920 -263 -880
rect -259 -920 -258 -880
rect -256 -920 -255 -880
rect -229 -887 -228 -847
rect -226 -887 -225 -847
rect -221 -887 -220 -847
rect -218 -887 -217 -847
rect -199 -858 -198 -838
rect -196 -858 -195 -838
rect 1349 -784 1350 -744
rect 1352 -784 1353 -744
rect 1357 -784 1358 -744
rect 1360 -784 1361 -744
rect 1387 -751 1388 -711
rect 1390 -751 1391 -711
rect 1395 -751 1396 -711
rect 1398 -751 1399 -711
rect 1417 -722 1418 -702
rect 1420 -722 1421 -702
rect 1514 -707 1515 -703
rect 1517 -707 1518 -703
rect 296 -792 297 -788
rect 299 -792 300 -788
rect -110 -917 -109 -897
rect -107 -917 -106 -897
rect -72 -940 -71 -900
rect -69 -940 -68 -900
rect -64 -940 -63 -900
rect -61 -940 -60 -900
rect -34 -907 -33 -867
rect -31 -907 -30 -867
rect -26 -907 -25 -867
rect -23 -907 -22 -867
rect -4 -878 -3 -858
rect -1 -878 0 -858
rect 230 -884 231 -880
rect 233 -884 234 -880
rect 246 -884 247 -880
rect 249 -884 257 -880
rect 259 -884 261 -880
rect 265 -884 267 -880
rect 269 -884 277 -880
rect 279 -884 280 -880
rect 296 -884 297 -880
rect 299 -884 300 -880
rect 527 -901 528 -897
rect 530 -901 538 -897
rect 540 -901 542 -897
rect 570 -901 571 -897
rect 573 -901 574 -897
rect 918 -899 919 -895
rect 921 -899 929 -895
rect 931 -899 939 -895
rect 941 -899 949 -895
rect 951 -899 959 -895
rect 961 -899 963 -895
rect 991 -899 992 -895
rect 994 -899 995 -895
rect 718 -933 719 -929
rect 721 -933 729 -929
rect 731 -933 739 -929
rect 741 -933 749 -929
rect 751 -933 753 -929
rect 779 -933 780 -929
rect 782 -933 783 -929
rect -307 -1088 -306 -1068
rect -304 -1088 -303 -1068
rect -269 -1111 -268 -1071
rect -266 -1111 -265 -1071
rect -261 -1111 -260 -1071
rect -258 -1111 -257 -1071
rect -231 -1078 -230 -1038
rect -228 -1078 -227 -1038
rect -223 -1078 -222 -1038
rect -220 -1078 -219 -1038
rect -201 -1049 -200 -1029
rect -198 -1049 -197 -1029
rect 230 -976 231 -972
rect 233 -976 234 -972
rect 246 -976 247 -972
rect 249 -976 257 -972
rect 259 -976 261 -972
rect 265 -976 267 -972
rect 269 -976 277 -972
rect 279 -976 280 -972
rect 296 -976 297 -972
rect 299 -976 300 -972
rect 1101 -960 1102 -956
rect 1104 -960 1105 -956
rect 1117 -960 1118 -956
rect 1120 -960 1128 -956
rect 1130 -960 1132 -956
rect 1136 -960 1138 -956
rect 1140 -960 1148 -956
rect 1150 -960 1151 -956
rect 1314 -951 1315 -931
rect 1317 -951 1318 -931
rect 1167 -960 1168 -956
rect 1170 -960 1171 -956
rect 1352 -974 1353 -934
rect 1355 -974 1356 -934
rect 1360 -974 1361 -934
rect 1363 -974 1364 -934
rect 1390 -941 1391 -901
rect 1393 -941 1394 -901
rect 1398 -941 1399 -901
rect 1401 -941 1402 -901
rect 1420 -912 1421 -892
rect 1423 -912 1424 -892
rect 1514 -897 1515 -893
rect 1517 -897 1518 -893
rect 526 -1006 527 -1002
rect 529 -1006 531 -1002
rect 535 -1006 537 -1002
rect 539 -1006 540 -1002
rect 554 -1006 555 -1002
rect 557 -1006 558 -1002
rect -109 -1100 -108 -1080
rect -106 -1100 -105 -1080
rect -71 -1123 -70 -1083
rect -68 -1123 -67 -1083
rect -63 -1123 -62 -1083
rect -60 -1123 -59 -1083
rect -33 -1090 -32 -1050
rect -30 -1090 -29 -1050
rect -25 -1090 -24 -1050
rect -22 -1090 -21 -1050
rect -3 -1061 -2 -1041
rect 0 -1061 1 -1041
rect 918 -998 919 -994
rect 921 -998 929 -994
rect 931 -998 939 -994
rect 941 -998 949 -994
rect 951 -998 953 -994
rect 979 -998 980 -994
rect 982 -998 983 -994
rect 718 -1030 719 -1026
rect 721 -1030 729 -1026
rect 731 -1030 739 -1026
rect 741 -1030 743 -1026
rect 771 -1030 772 -1026
rect 774 -1030 775 -1026
rect 230 -1069 231 -1065
rect 233 -1069 234 -1065
rect 246 -1069 247 -1065
rect 249 -1069 257 -1065
rect 259 -1069 261 -1065
rect 265 -1069 267 -1065
rect 269 -1069 277 -1065
rect 279 -1069 280 -1065
rect 296 -1069 297 -1065
rect 299 -1069 300 -1065
rect 1101 -1058 1102 -1054
rect 1104 -1058 1105 -1054
rect 1117 -1058 1118 -1054
rect 1120 -1058 1128 -1054
rect 1130 -1058 1132 -1054
rect 1136 -1058 1138 -1054
rect 1140 -1058 1148 -1054
rect 1150 -1058 1151 -1054
rect 531 -1089 532 -1085
rect 534 -1089 542 -1085
rect 544 -1089 552 -1085
rect 554 -1089 556 -1085
rect 584 -1089 585 -1085
rect 587 -1089 588 -1085
rect 1167 -1058 1168 -1054
rect 1170 -1058 1171 -1054
rect 918 -1091 919 -1087
rect 921 -1091 929 -1087
rect 931 -1091 939 -1087
rect 941 -1091 943 -1087
rect 971 -1091 972 -1087
rect 974 -1091 975 -1087
rect 717 -1118 718 -1114
rect 720 -1118 728 -1114
rect 730 -1118 732 -1114
rect 760 -1118 761 -1114
rect 763 -1118 764 -1114
rect 240 -1157 241 -1153
rect 243 -1157 251 -1153
rect 253 -1157 255 -1153
rect 283 -1157 284 -1153
rect 286 -1157 287 -1153
rect -307 -1282 -306 -1262
rect -304 -1282 -303 -1262
rect -269 -1305 -268 -1265
rect -266 -1305 -265 -1265
rect -261 -1305 -260 -1265
rect -258 -1305 -257 -1265
rect -231 -1272 -230 -1232
rect -228 -1272 -227 -1232
rect -223 -1272 -222 -1232
rect -220 -1272 -219 -1232
rect -201 -1243 -200 -1223
rect -198 -1243 -197 -1223
rect 531 -1172 532 -1168
rect 534 -1172 542 -1168
rect 544 -1172 546 -1168
rect 574 -1172 575 -1168
rect 577 -1172 578 -1168
rect -105 -1282 -104 -1262
rect -102 -1282 -101 -1262
rect -67 -1305 -66 -1265
rect -64 -1305 -63 -1265
rect -59 -1305 -58 -1265
rect -56 -1305 -55 -1265
rect -29 -1272 -28 -1232
rect -26 -1272 -25 -1232
rect -21 -1272 -20 -1232
rect -18 -1272 -17 -1232
rect 1 -1243 2 -1223
rect 4 -1243 5 -1223
rect 1312 -1140 1313 -1120
rect 1315 -1140 1316 -1120
rect 1101 -1158 1102 -1154
rect 1104 -1158 1105 -1154
rect 1117 -1158 1118 -1154
rect 1120 -1158 1128 -1154
rect 1130 -1158 1132 -1154
rect 1136 -1158 1138 -1154
rect 1140 -1158 1148 -1154
rect 1150 -1158 1151 -1154
rect 1167 -1158 1168 -1154
rect 1170 -1158 1171 -1154
rect 1350 -1163 1351 -1123
rect 1353 -1163 1354 -1123
rect 1358 -1163 1359 -1123
rect 1361 -1163 1362 -1123
rect 1388 -1130 1389 -1090
rect 1391 -1130 1392 -1090
rect 1396 -1130 1397 -1090
rect 1399 -1130 1400 -1090
rect 1418 -1101 1419 -1081
rect 1421 -1101 1422 -1081
rect 1513 -1086 1514 -1082
rect 1516 -1086 1517 -1082
rect 916 -1175 917 -1171
rect 919 -1175 927 -1171
rect 929 -1175 931 -1171
rect 959 -1175 960 -1171
rect 962 -1175 963 -1171
rect 715 -1217 716 -1213
rect 718 -1217 720 -1213
rect 724 -1217 726 -1213
rect 728 -1217 729 -1213
rect 733 -1217 735 -1213
rect 737 -1217 739 -1213
rect 743 -1217 745 -1213
rect 747 -1217 749 -1213
rect 763 -1217 764 -1213
rect 766 -1217 767 -1213
rect 239 -1232 240 -1228
rect 242 -1232 250 -1228
rect 252 -1232 254 -1228
rect 282 -1232 283 -1228
rect 285 -1232 286 -1228
rect 530 -1264 531 -1260
rect 533 -1264 535 -1260
rect 539 -1264 541 -1260
rect 543 -1264 544 -1260
rect 548 -1264 550 -1260
rect 552 -1264 554 -1260
rect 568 -1264 569 -1260
rect 571 -1264 572 -1260
rect 1101 -1256 1102 -1252
rect 1104 -1256 1105 -1252
rect 1117 -1256 1118 -1252
rect 1120 -1256 1128 -1252
rect 1130 -1256 1132 -1252
rect 1136 -1256 1138 -1252
rect 1140 -1256 1148 -1252
rect 1150 -1256 1151 -1252
rect 1167 -1256 1168 -1252
rect 1170 -1256 1171 -1252
rect 915 -1293 916 -1289
rect 918 -1293 920 -1289
rect 924 -1293 926 -1289
rect 928 -1293 929 -1289
rect 933 -1293 935 -1289
rect 937 -1293 939 -1289
rect 943 -1293 945 -1289
rect 947 -1293 949 -1289
rect 953 -1293 955 -1289
rect 957 -1293 959 -1289
rect 972 -1293 973 -1289
rect 975 -1293 976 -1289
rect 239 -1307 240 -1303
rect 242 -1307 250 -1303
rect 252 -1307 254 -1303
rect 282 -1307 283 -1303
rect 285 -1307 286 -1303
rect 1313 -1329 1314 -1309
rect 1316 -1329 1317 -1309
rect -307 -1466 -306 -1446
rect -304 -1466 -303 -1446
rect -269 -1489 -268 -1449
rect -266 -1489 -265 -1449
rect -261 -1489 -260 -1449
rect -258 -1489 -257 -1449
rect -231 -1456 -230 -1416
rect -228 -1456 -227 -1416
rect -223 -1456 -222 -1416
rect -220 -1456 -219 -1416
rect -201 -1427 -200 -1407
rect -198 -1427 -197 -1407
rect 1351 -1352 1352 -1312
rect 1354 -1352 1355 -1312
rect 1359 -1352 1360 -1312
rect 1362 -1352 1363 -1312
rect 1389 -1319 1390 -1279
rect 1392 -1319 1393 -1279
rect 1397 -1319 1398 -1279
rect 1400 -1319 1401 -1279
rect 1419 -1290 1420 -1270
rect 1422 -1290 1423 -1270
rect 1511 -1275 1512 -1271
rect 1514 -1275 1515 -1271
rect 239 -1382 240 -1378
rect 242 -1382 250 -1378
rect 252 -1382 254 -1378
rect 282 -1382 283 -1378
rect 285 -1382 286 -1378
rect -102 -1464 -101 -1444
rect -99 -1464 -98 -1444
rect -64 -1487 -63 -1447
rect -61 -1487 -60 -1447
rect -56 -1487 -55 -1447
rect -53 -1487 -52 -1447
rect -26 -1454 -25 -1414
rect -23 -1454 -22 -1414
rect -18 -1454 -17 -1414
rect -15 -1454 -14 -1414
rect 4 -1425 5 -1405
rect 7 -1425 8 -1405
rect 1314 -1517 1315 -1497
rect 1317 -1517 1318 -1497
rect 1352 -1540 1353 -1500
rect 1355 -1540 1356 -1500
rect 1360 -1540 1361 -1500
rect 1363 -1540 1364 -1500
rect 1390 -1507 1391 -1467
rect 1393 -1507 1394 -1467
rect 1398 -1507 1399 -1467
rect 1401 -1507 1402 -1467
rect 1420 -1478 1421 -1458
rect 1423 -1478 1424 -1458
rect 1514 -1463 1515 -1459
rect 1517 -1463 1518 -1459
<< pdiffusion >>
rect 1311 -726 1312 -646
rect 1314 -726 1315 -646
rect 1319 -726 1320 -646
rect 1322 -726 1323 -646
rect 1349 -726 1350 -646
rect 1352 -726 1353 -646
rect 1357 -726 1358 -646
rect 1360 -726 1361 -646
rect 1387 -696 1388 -646
rect 1390 -696 1391 -646
rect 1417 -688 1418 -648
rect 1420 -688 1421 -648
rect 1514 -688 1515 -680
rect 1517 -688 1518 -680
rect 230 -746 231 -740
rect 233 -746 234 -740
rect 246 -746 247 -740
rect 249 -746 257 -740
rect 259 -746 261 -740
rect 265 -746 267 -740
rect 269 -746 277 -740
rect 279 -746 280 -740
rect 296 -746 297 -740
rect 299 -746 300 -740
rect -305 -862 -304 -782
rect -302 -862 -301 -782
rect -297 -862 -296 -782
rect -294 -862 -293 -782
rect -267 -862 -266 -782
rect -264 -862 -263 -782
rect -259 -862 -258 -782
rect -256 -862 -255 -782
rect -229 -832 -228 -782
rect -226 -832 -225 -782
rect -199 -824 -198 -784
rect -196 -824 -195 -784
rect -110 -882 -109 -802
rect -107 -882 -106 -802
rect -102 -882 -101 -802
rect -99 -882 -98 -802
rect -72 -882 -71 -802
rect -69 -882 -68 -802
rect -64 -882 -63 -802
rect -61 -882 -60 -802
rect -34 -852 -33 -802
rect -31 -852 -30 -802
rect -4 -844 -3 -804
rect -1 -844 0 -804
rect 230 -838 231 -832
rect 233 -838 234 -832
rect 246 -838 247 -832
rect 249 -838 257 -832
rect 259 -838 261 -832
rect 265 -838 267 -832
rect 269 -838 277 -832
rect 279 -838 280 -832
rect 296 -838 297 -832
rect 299 -838 300 -832
rect 918 -851 919 -845
rect 921 -851 923 -845
rect 927 -851 929 -845
rect 931 -851 933 -845
rect 937 -851 939 -845
rect 941 -851 943 -845
rect 947 -851 949 -845
rect 951 -851 953 -845
rect 957 -851 959 -845
rect 961 -851 963 -845
rect 991 -851 992 -845
rect 994 -851 995 -845
rect 527 -871 528 -865
rect 530 -871 532 -865
rect 536 -871 538 -865
rect 540 -871 542 -865
rect 570 -871 571 -865
rect 573 -871 574 -865
rect 718 -892 719 -886
rect 721 -892 723 -886
rect 727 -892 729 -886
rect 731 -892 733 -886
rect 737 -892 739 -886
rect 741 -892 743 -886
rect 747 -892 749 -886
rect 751 -892 753 -886
rect 779 -892 780 -886
rect 782 -892 783 -886
rect 230 -930 231 -924
rect 233 -930 234 -924
rect 246 -930 247 -924
rect 249 -930 257 -924
rect 259 -930 261 -924
rect 265 -930 267 -924
rect 269 -930 277 -924
rect 279 -930 280 -924
rect 296 -930 297 -924
rect 299 -930 300 -924
rect -307 -1053 -306 -973
rect -304 -1053 -303 -973
rect -299 -1053 -298 -973
rect -296 -1053 -295 -973
rect -269 -1053 -268 -973
rect -266 -1053 -265 -973
rect -261 -1053 -260 -973
rect -258 -1053 -257 -973
rect -231 -1023 -230 -973
rect -228 -1023 -227 -973
rect 1101 -914 1102 -908
rect 1104 -914 1105 -908
rect 1117 -914 1118 -908
rect 1120 -914 1128 -908
rect 1130 -914 1132 -908
rect 1136 -914 1138 -908
rect 1140 -914 1148 -908
rect 1150 -914 1151 -908
rect 1167 -914 1168 -908
rect 1170 -914 1171 -908
rect 918 -957 919 -951
rect 921 -957 923 -951
rect 927 -957 929 -951
rect 931 -957 933 -951
rect 937 -957 939 -951
rect 941 -957 943 -951
rect 947 -957 949 -951
rect 951 -957 953 -951
rect 979 -957 980 -951
rect 982 -957 983 -951
rect 1314 -916 1315 -836
rect 1317 -916 1318 -836
rect 1322 -916 1323 -836
rect 1325 -916 1326 -836
rect 1352 -916 1353 -836
rect 1355 -916 1356 -836
rect 1360 -916 1361 -836
rect 1363 -916 1364 -836
rect 1390 -886 1391 -836
rect 1393 -886 1394 -836
rect 1420 -878 1421 -838
rect 1423 -878 1424 -838
rect 1514 -878 1515 -870
rect 1517 -878 1518 -870
rect -201 -1015 -200 -975
rect -198 -1015 -197 -975
rect -109 -1065 -108 -985
rect -106 -1065 -105 -985
rect -101 -1065 -100 -985
rect -98 -1065 -97 -985
rect -71 -1065 -70 -985
rect -68 -1065 -67 -985
rect -63 -1065 -62 -985
rect -60 -1065 -59 -985
rect -33 -1035 -32 -985
rect -30 -1035 -29 -985
rect 526 -970 527 -964
rect 529 -970 537 -964
rect 539 -970 540 -964
rect 554 -970 555 -964
rect 557 -970 558 -964
rect -3 -1027 -2 -987
rect 0 -1027 1 -987
rect 718 -997 719 -991
rect 721 -997 723 -991
rect 727 -997 729 -991
rect 731 -997 733 -991
rect 737 -997 739 -991
rect 741 -997 743 -991
rect 771 -997 772 -991
rect 774 -997 775 -991
rect 230 -1023 231 -1017
rect 233 -1023 234 -1017
rect 246 -1023 247 -1017
rect 249 -1023 257 -1017
rect 259 -1023 261 -1017
rect 265 -1023 267 -1017
rect 269 -1023 277 -1017
rect 279 -1023 280 -1017
rect 296 -1023 297 -1017
rect 299 -1023 300 -1017
rect 1101 -1012 1102 -1006
rect 1104 -1012 1105 -1006
rect 1117 -1012 1118 -1006
rect 1120 -1012 1128 -1006
rect 1130 -1012 1132 -1006
rect 1136 -1012 1138 -1006
rect 1140 -1012 1148 -1006
rect 1150 -1012 1151 -1006
rect 1167 -1012 1168 -1006
rect 1170 -1012 1171 -1006
rect 531 -1056 532 -1050
rect 534 -1056 536 -1050
rect 540 -1056 542 -1050
rect 544 -1056 546 -1050
rect 550 -1056 552 -1050
rect 554 -1056 556 -1050
rect 584 -1056 585 -1050
rect 587 -1056 588 -1050
rect 918 -1058 919 -1052
rect 921 -1058 923 -1052
rect 927 -1058 929 -1052
rect 931 -1058 933 -1052
rect 937 -1058 939 -1052
rect 941 -1058 943 -1052
rect 971 -1058 972 -1052
rect 974 -1058 975 -1052
rect 717 -1088 718 -1082
rect 720 -1088 722 -1082
rect 726 -1088 728 -1082
rect 730 -1088 732 -1082
rect 760 -1088 761 -1082
rect 763 -1088 764 -1082
rect 1101 -1112 1102 -1106
rect 1104 -1112 1105 -1106
rect 1117 -1112 1118 -1106
rect 1120 -1112 1128 -1106
rect 1130 -1112 1132 -1106
rect 1136 -1112 1138 -1106
rect 1140 -1112 1148 -1106
rect 1150 -1112 1151 -1106
rect 1167 -1112 1168 -1106
rect 1170 -1112 1171 -1106
rect 240 -1127 241 -1121
rect 243 -1127 245 -1121
rect 249 -1127 251 -1121
rect 253 -1127 255 -1121
rect 283 -1127 284 -1121
rect 286 -1127 287 -1121
rect 531 -1142 532 -1136
rect 534 -1142 536 -1136
rect 540 -1142 542 -1136
rect 544 -1142 546 -1136
rect 574 -1142 575 -1136
rect 577 -1142 578 -1136
rect -307 -1247 -306 -1167
rect -304 -1247 -303 -1167
rect -299 -1247 -298 -1167
rect -296 -1247 -295 -1167
rect -269 -1247 -268 -1167
rect -266 -1247 -265 -1167
rect -261 -1247 -260 -1167
rect -258 -1247 -257 -1167
rect -231 -1217 -230 -1167
rect -228 -1217 -227 -1167
rect -201 -1209 -200 -1169
rect -198 -1209 -197 -1169
rect -105 -1247 -104 -1167
rect -102 -1247 -101 -1167
rect -97 -1247 -96 -1167
rect -94 -1247 -93 -1167
rect -67 -1247 -66 -1167
rect -64 -1247 -63 -1167
rect -59 -1247 -58 -1167
rect -56 -1247 -55 -1167
rect -29 -1217 -28 -1167
rect -26 -1217 -25 -1167
rect 916 -1145 917 -1139
rect 919 -1145 921 -1139
rect 925 -1145 927 -1139
rect 929 -1145 931 -1139
rect 959 -1145 960 -1139
rect 962 -1145 963 -1139
rect 715 -1167 716 -1161
rect 718 -1167 726 -1161
rect 728 -1167 735 -1161
rect 737 -1167 745 -1161
rect 747 -1167 749 -1161
rect 763 -1167 764 -1161
rect 766 -1167 767 -1161
rect 1 -1209 2 -1169
rect 4 -1209 5 -1169
rect 239 -1202 240 -1196
rect 242 -1202 244 -1196
rect 248 -1202 250 -1196
rect 252 -1202 254 -1196
rect 282 -1202 283 -1196
rect 285 -1202 286 -1196
rect 1312 -1105 1313 -1025
rect 1315 -1105 1316 -1025
rect 1320 -1105 1321 -1025
rect 1323 -1105 1324 -1025
rect 1350 -1105 1351 -1025
rect 1353 -1105 1354 -1025
rect 1358 -1105 1359 -1025
rect 1361 -1105 1362 -1025
rect 1388 -1075 1389 -1025
rect 1391 -1075 1392 -1025
rect 1418 -1067 1419 -1027
rect 1421 -1067 1422 -1027
rect 1513 -1067 1514 -1059
rect 1516 -1067 1517 -1059
rect 1101 -1210 1102 -1204
rect 1104 -1210 1105 -1204
rect 1117 -1210 1118 -1204
rect 1120 -1210 1128 -1204
rect 1130 -1210 1132 -1204
rect 1136 -1210 1138 -1204
rect 1140 -1210 1148 -1204
rect 1150 -1210 1151 -1204
rect 1167 -1210 1168 -1204
rect 1170 -1210 1171 -1204
rect 530 -1221 531 -1215
rect 533 -1221 541 -1215
rect 543 -1221 550 -1215
rect 552 -1221 554 -1215
rect 568 -1221 569 -1215
rect 571 -1221 572 -1215
rect 915 -1236 916 -1230
rect 918 -1236 926 -1230
rect 928 -1236 935 -1230
rect 937 -1236 945 -1230
rect 947 -1236 955 -1230
rect 957 -1236 959 -1230
rect 972 -1236 973 -1230
rect 975 -1236 976 -1230
rect 239 -1277 240 -1271
rect 242 -1277 244 -1271
rect 248 -1277 250 -1271
rect 252 -1277 254 -1271
rect 282 -1277 283 -1271
rect 285 -1277 286 -1271
rect 1313 -1294 1314 -1214
rect 1316 -1294 1317 -1214
rect 1321 -1294 1322 -1214
rect 1324 -1294 1325 -1214
rect 1351 -1294 1352 -1214
rect 1354 -1294 1355 -1214
rect 1359 -1294 1360 -1214
rect 1362 -1294 1363 -1214
rect 1389 -1264 1390 -1214
rect 1392 -1264 1393 -1214
rect 1419 -1256 1420 -1216
rect 1422 -1256 1423 -1216
rect 1511 -1256 1512 -1248
rect 1514 -1256 1515 -1248
rect -307 -1431 -306 -1351
rect -304 -1431 -303 -1351
rect -299 -1431 -298 -1351
rect -296 -1431 -295 -1351
rect -269 -1431 -268 -1351
rect -266 -1431 -265 -1351
rect -261 -1431 -260 -1351
rect -258 -1431 -257 -1351
rect -231 -1401 -230 -1351
rect -228 -1401 -227 -1351
rect -201 -1393 -200 -1353
rect -198 -1393 -197 -1353
rect -102 -1429 -101 -1349
rect -99 -1429 -98 -1349
rect -94 -1429 -93 -1349
rect -91 -1429 -90 -1349
rect -64 -1429 -63 -1349
rect -61 -1429 -60 -1349
rect -56 -1429 -55 -1349
rect -53 -1429 -52 -1349
rect -26 -1399 -25 -1349
rect -23 -1399 -22 -1349
rect 4 -1391 5 -1351
rect 7 -1391 8 -1351
rect 239 -1352 240 -1346
rect 242 -1352 244 -1346
rect 248 -1352 250 -1346
rect 252 -1352 254 -1346
rect 282 -1352 283 -1346
rect 285 -1352 286 -1346
rect 1314 -1482 1315 -1402
rect 1317 -1482 1318 -1402
rect 1322 -1482 1323 -1402
rect 1325 -1482 1326 -1402
rect 1352 -1482 1353 -1402
rect 1355 -1482 1356 -1402
rect 1360 -1482 1361 -1402
rect 1363 -1482 1364 -1402
rect 1390 -1452 1391 -1402
rect 1393 -1452 1394 -1402
rect 1420 -1444 1421 -1404
rect 1423 -1444 1424 -1404
rect 1514 -1444 1515 -1436
rect 1517 -1444 1518 -1436
<< ndcontact >>
rect 1307 -761 1311 -741
rect 1315 -761 1319 -741
rect 226 -792 230 -788
rect 234 -792 238 -788
rect 242 -792 246 -788
rect 261 -792 265 -788
rect 280 -792 284 -788
rect -309 -897 -305 -877
rect -301 -897 -297 -877
rect -271 -920 -267 -880
rect -263 -920 -259 -880
rect -255 -920 -251 -880
rect -233 -887 -229 -847
rect -225 -887 -221 -847
rect -217 -887 -213 -847
rect -203 -858 -199 -838
rect -195 -858 -191 -838
rect 1345 -784 1349 -744
rect 1353 -784 1357 -744
rect 1361 -784 1365 -744
rect 1383 -751 1387 -711
rect 1391 -751 1395 -711
rect 1399 -751 1403 -711
rect 1413 -722 1417 -702
rect 1421 -722 1425 -702
rect 1510 -707 1514 -703
rect 1518 -707 1522 -703
rect 292 -792 296 -788
rect 300 -792 304 -788
rect -114 -917 -110 -897
rect -106 -917 -102 -897
rect -76 -940 -72 -900
rect -68 -940 -64 -900
rect -60 -940 -56 -900
rect -38 -907 -34 -867
rect -30 -907 -26 -867
rect -22 -907 -18 -867
rect -8 -878 -4 -858
rect 0 -878 4 -858
rect 226 -884 230 -880
rect 234 -884 238 -880
rect 242 -884 246 -880
rect 261 -884 265 -880
rect 280 -884 284 -880
rect 292 -884 296 -880
rect 300 -884 304 -880
rect 523 -901 527 -897
rect 542 -901 546 -897
rect 566 -901 570 -897
rect 574 -901 578 -897
rect 914 -899 918 -895
rect 963 -899 967 -895
rect 987 -899 991 -895
rect 995 -899 999 -895
rect 714 -933 718 -929
rect 753 -933 757 -929
rect 775 -933 779 -929
rect 783 -933 787 -929
rect -311 -1088 -307 -1068
rect -303 -1088 -299 -1068
rect -273 -1111 -269 -1071
rect -265 -1111 -261 -1071
rect -257 -1111 -253 -1071
rect -235 -1078 -231 -1038
rect -227 -1078 -223 -1038
rect -219 -1078 -215 -1038
rect -205 -1049 -201 -1029
rect -197 -1049 -193 -1029
rect 226 -976 230 -972
rect 234 -976 238 -972
rect 242 -976 246 -972
rect 261 -976 265 -972
rect 280 -976 284 -972
rect 292 -976 296 -972
rect 300 -976 304 -972
rect 1097 -960 1101 -956
rect 1105 -960 1109 -956
rect 1113 -960 1117 -956
rect 1132 -960 1136 -956
rect 1151 -960 1155 -956
rect 1310 -951 1314 -931
rect 1318 -951 1322 -931
rect 1163 -960 1167 -956
rect 1171 -960 1175 -956
rect 1348 -974 1352 -934
rect 1356 -974 1360 -934
rect 1364 -974 1368 -934
rect 1386 -941 1390 -901
rect 1394 -941 1398 -901
rect 1402 -941 1406 -901
rect 1416 -912 1420 -892
rect 1424 -912 1428 -892
rect 1510 -897 1514 -893
rect 1518 -897 1522 -893
rect 522 -1006 526 -1002
rect 531 -1006 535 -1002
rect 540 -1006 544 -1002
rect 550 -1006 554 -1002
rect 558 -1006 562 -1002
rect -113 -1100 -109 -1080
rect -105 -1100 -101 -1080
rect -75 -1123 -71 -1083
rect -67 -1123 -63 -1083
rect -59 -1123 -55 -1083
rect -37 -1090 -33 -1050
rect -29 -1090 -25 -1050
rect -21 -1090 -17 -1050
rect -7 -1061 -3 -1041
rect 1 -1061 5 -1041
rect 914 -998 918 -994
rect 953 -998 957 -994
rect 975 -998 979 -994
rect 983 -998 987 -994
rect 714 -1030 718 -1026
rect 743 -1030 747 -1026
rect 767 -1030 771 -1026
rect 775 -1030 779 -1026
rect 226 -1069 230 -1065
rect 234 -1069 238 -1065
rect 242 -1069 246 -1065
rect 261 -1069 265 -1065
rect 280 -1069 284 -1065
rect 292 -1069 296 -1065
rect 300 -1069 304 -1065
rect 1097 -1058 1101 -1054
rect 1105 -1058 1109 -1054
rect 1113 -1058 1117 -1054
rect 1132 -1058 1136 -1054
rect 1151 -1058 1155 -1054
rect 527 -1089 531 -1085
rect 556 -1089 560 -1085
rect 580 -1089 584 -1085
rect 588 -1089 592 -1085
rect 1163 -1058 1167 -1054
rect 1171 -1058 1175 -1054
rect 914 -1091 918 -1087
rect 943 -1091 947 -1087
rect 967 -1091 971 -1087
rect 975 -1091 979 -1087
rect 713 -1118 717 -1114
rect 732 -1118 736 -1114
rect 756 -1118 760 -1114
rect 764 -1118 768 -1114
rect 236 -1157 240 -1153
rect 255 -1157 259 -1153
rect 279 -1157 283 -1153
rect 287 -1157 291 -1153
rect -311 -1282 -307 -1262
rect -303 -1282 -299 -1262
rect -273 -1305 -269 -1265
rect -265 -1305 -261 -1265
rect -257 -1305 -253 -1265
rect -235 -1272 -231 -1232
rect -227 -1272 -223 -1232
rect -219 -1272 -215 -1232
rect -205 -1243 -201 -1223
rect -197 -1243 -193 -1223
rect 527 -1172 531 -1168
rect 546 -1172 550 -1168
rect 570 -1172 574 -1168
rect 578 -1172 582 -1168
rect -109 -1282 -105 -1262
rect -101 -1282 -97 -1262
rect -71 -1305 -67 -1265
rect -63 -1305 -59 -1265
rect -55 -1305 -51 -1265
rect -33 -1272 -29 -1232
rect -25 -1272 -21 -1232
rect -17 -1272 -13 -1232
rect -3 -1243 1 -1223
rect 5 -1243 9 -1223
rect 1308 -1140 1312 -1120
rect 1316 -1140 1320 -1120
rect 1097 -1158 1101 -1154
rect 1105 -1158 1109 -1154
rect 1113 -1158 1117 -1154
rect 1132 -1158 1136 -1154
rect 1151 -1158 1155 -1154
rect 1163 -1158 1167 -1154
rect 1171 -1158 1175 -1154
rect 1346 -1163 1350 -1123
rect 1354 -1163 1358 -1123
rect 1362 -1163 1366 -1123
rect 1384 -1130 1388 -1090
rect 1392 -1130 1396 -1090
rect 1400 -1130 1404 -1090
rect 1414 -1101 1418 -1081
rect 1422 -1101 1426 -1081
rect 1509 -1086 1513 -1082
rect 1517 -1086 1521 -1082
rect 912 -1175 916 -1171
rect 931 -1175 935 -1171
rect 955 -1175 959 -1171
rect 963 -1175 967 -1171
rect 711 -1217 715 -1213
rect 720 -1217 724 -1213
rect 729 -1217 733 -1213
rect 739 -1217 743 -1213
rect 749 -1217 753 -1213
rect 759 -1217 763 -1213
rect 767 -1217 771 -1213
rect 235 -1232 239 -1228
rect 254 -1232 258 -1228
rect 278 -1232 282 -1228
rect 286 -1232 290 -1228
rect 526 -1264 530 -1260
rect 535 -1264 539 -1260
rect 544 -1264 548 -1260
rect 554 -1264 558 -1260
rect 564 -1264 568 -1260
rect 572 -1264 576 -1260
rect 1097 -1256 1101 -1252
rect 1105 -1256 1109 -1252
rect 1113 -1256 1117 -1252
rect 1132 -1256 1136 -1252
rect 1151 -1256 1155 -1252
rect 1163 -1256 1167 -1252
rect 1171 -1256 1175 -1252
rect 911 -1293 915 -1289
rect 920 -1293 924 -1289
rect 929 -1293 933 -1289
rect 939 -1293 943 -1289
rect 949 -1293 953 -1289
rect 959 -1293 963 -1289
rect 968 -1293 972 -1289
rect 976 -1293 980 -1289
rect 235 -1307 239 -1303
rect 254 -1307 258 -1303
rect 278 -1307 282 -1303
rect 286 -1307 290 -1303
rect 1309 -1329 1313 -1309
rect 1317 -1329 1321 -1309
rect -311 -1466 -307 -1446
rect -303 -1466 -299 -1446
rect -273 -1489 -269 -1449
rect -265 -1489 -261 -1449
rect -257 -1489 -253 -1449
rect -235 -1456 -231 -1416
rect -227 -1456 -223 -1416
rect -219 -1456 -215 -1416
rect -205 -1427 -201 -1407
rect -197 -1427 -193 -1407
rect 1347 -1352 1351 -1312
rect 1355 -1352 1359 -1312
rect 1363 -1352 1367 -1312
rect 1385 -1319 1389 -1279
rect 1393 -1319 1397 -1279
rect 1401 -1319 1405 -1279
rect 1415 -1290 1419 -1270
rect 1423 -1290 1427 -1270
rect 1507 -1275 1511 -1271
rect 1515 -1275 1519 -1271
rect 235 -1382 239 -1378
rect 254 -1382 258 -1378
rect 278 -1382 282 -1378
rect 286 -1382 290 -1378
rect -106 -1464 -102 -1444
rect -98 -1464 -94 -1444
rect -68 -1487 -64 -1447
rect -60 -1487 -56 -1447
rect -52 -1487 -48 -1447
rect -30 -1454 -26 -1414
rect -22 -1454 -18 -1414
rect -14 -1454 -10 -1414
rect 0 -1425 4 -1405
rect 8 -1425 12 -1405
rect 1310 -1517 1314 -1497
rect 1318 -1517 1322 -1497
rect 1348 -1540 1352 -1500
rect 1356 -1540 1360 -1500
rect 1364 -1540 1368 -1500
rect 1386 -1507 1390 -1467
rect 1394 -1507 1398 -1467
rect 1402 -1507 1406 -1467
rect 1416 -1478 1420 -1458
rect 1424 -1478 1428 -1458
rect 1510 -1463 1514 -1459
rect 1518 -1463 1522 -1459
<< pdcontact >>
rect 1307 -726 1311 -646
rect 1315 -726 1319 -646
rect 1323 -726 1327 -646
rect 1345 -726 1349 -646
rect 1353 -726 1357 -646
rect 1361 -726 1365 -646
rect 1383 -696 1387 -646
rect 1391 -696 1395 -646
rect 1413 -688 1417 -648
rect 1421 -688 1425 -648
rect 1510 -688 1514 -680
rect 1518 -688 1522 -680
rect 226 -746 230 -740
rect 234 -746 238 -740
rect 242 -746 246 -740
rect 261 -746 265 -740
rect 280 -746 284 -740
rect 292 -746 296 -740
rect 300 -746 304 -740
rect -309 -862 -305 -782
rect -301 -862 -297 -782
rect -293 -862 -289 -782
rect -271 -862 -267 -782
rect -263 -862 -259 -782
rect -255 -862 -251 -782
rect -233 -832 -229 -782
rect -225 -832 -221 -782
rect -203 -824 -199 -784
rect -195 -824 -191 -784
rect -114 -882 -110 -802
rect -106 -882 -102 -802
rect -98 -882 -94 -802
rect -76 -882 -72 -802
rect -68 -882 -64 -802
rect -60 -882 -56 -802
rect -38 -852 -34 -802
rect -30 -852 -26 -802
rect -8 -844 -4 -804
rect 0 -844 4 -804
rect 226 -838 230 -832
rect 234 -838 238 -832
rect 242 -838 246 -832
rect 261 -838 265 -832
rect 280 -838 284 -832
rect 292 -838 296 -832
rect 300 -838 304 -832
rect 914 -851 918 -845
rect 923 -851 927 -845
rect 933 -851 937 -845
rect 943 -851 947 -845
rect 953 -851 957 -845
rect 963 -851 967 -845
rect 987 -851 991 -845
rect 995 -851 999 -845
rect 523 -871 527 -865
rect 532 -871 536 -865
rect 542 -871 546 -865
rect 566 -871 570 -865
rect 574 -871 578 -865
rect 714 -892 718 -886
rect 723 -892 727 -886
rect 733 -892 737 -886
rect 743 -892 747 -886
rect 753 -892 757 -886
rect 775 -892 779 -886
rect 783 -892 787 -886
rect 226 -930 230 -924
rect 234 -930 238 -924
rect 242 -930 246 -924
rect 261 -930 265 -924
rect 280 -930 284 -924
rect 292 -930 296 -924
rect 300 -930 304 -924
rect -311 -1053 -307 -973
rect -303 -1053 -299 -973
rect -295 -1053 -291 -973
rect -273 -1053 -269 -973
rect -265 -1053 -261 -973
rect -257 -1053 -253 -973
rect -235 -1023 -231 -973
rect -227 -1023 -223 -973
rect 1097 -914 1101 -908
rect 1105 -914 1109 -908
rect 1113 -914 1117 -908
rect 1132 -914 1136 -908
rect 1151 -914 1155 -908
rect 1163 -914 1167 -908
rect 1171 -914 1175 -908
rect 914 -957 918 -951
rect 923 -957 927 -951
rect 933 -957 937 -951
rect 943 -957 947 -951
rect 953 -957 957 -951
rect 975 -957 979 -951
rect 983 -957 987 -951
rect 1310 -916 1314 -836
rect 1318 -916 1322 -836
rect 1326 -916 1330 -836
rect 1348 -916 1352 -836
rect 1356 -916 1360 -836
rect 1364 -916 1368 -836
rect 1386 -886 1390 -836
rect 1394 -886 1398 -836
rect 1416 -878 1420 -838
rect 1424 -878 1428 -838
rect 1510 -878 1514 -870
rect 1518 -878 1522 -870
rect -205 -1015 -201 -975
rect -197 -1015 -193 -975
rect -113 -1065 -109 -985
rect -105 -1065 -101 -985
rect -97 -1065 -93 -985
rect -75 -1065 -71 -985
rect -67 -1065 -63 -985
rect -59 -1065 -55 -985
rect -37 -1035 -33 -985
rect -29 -1035 -25 -985
rect 522 -970 526 -964
rect 540 -970 544 -964
rect 550 -970 554 -964
rect 558 -970 562 -964
rect -7 -1027 -3 -987
rect 1 -1027 5 -987
rect 714 -997 718 -991
rect 723 -997 727 -991
rect 733 -997 737 -991
rect 743 -997 747 -991
rect 767 -997 771 -991
rect 775 -997 779 -991
rect 226 -1023 230 -1017
rect 234 -1023 238 -1017
rect 242 -1023 246 -1017
rect 261 -1023 265 -1017
rect 280 -1023 284 -1017
rect 292 -1023 296 -1017
rect 300 -1023 304 -1017
rect 1097 -1012 1101 -1006
rect 1105 -1012 1109 -1006
rect 1113 -1012 1117 -1006
rect 1132 -1012 1136 -1006
rect 1151 -1012 1155 -1006
rect 1163 -1012 1167 -1006
rect 1171 -1012 1175 -1006
rect 527 -1056 531 -1050
rect 536 -1056 540 -1050
rect 546 -1056 550 -1050
rect 556 -1056 560 -1050
rect 580 -1056 584 -1050
rect 588 -1056 592 -1050
rect 914 -1058 918 -1052
rect 923 -1058 927 -1052
rect 933 -1058 937 -1052
rect 943 -1058 947 -1052
rect 967 -1058 971 -1052
rect 975 -1058 979 -1052
rect 713 -1088 717 -1082
rect 722 -1088 726 -1082
rect 732 -1088 736 -1082
rect 756 -1088 760 -1082
rect 764 -1088 768 -1082
rect 1097 -1112 1101 -1106
rect 1105 -1112 1109 -1106
rect 1113 -1112 1117 -1106
rect 1132 -1112 1136 -1106
rect 1151 -1112 1155 -1106
rect 1163 -1112 1167 -1106
rect 1171 -1112 1175 -1106
rect 236 -1127 240 -1121
rect 245 -1127 249 -1121
rect 255 -1127 259 -1121
rect 279 -1127 283 -1121
rect 287 -1127 291 -1121
rect 527 -1142 531 -1136
rect 536 -1142 540 -1136
rect 546 -1142 550 -1136
rect 570 -1142 574 -1136
rect 578 -1142 582 -1136
rect -311 -1247 -307 -1167
rect -303 -1247 -299 -1167
rect -295 -1247 -291 -1167
rect -273 -1247 -269 -1167
rect -265 -1247 -261 -1167
rect -257 -1247 -253 -1167
rect -235 -1217 -231 -1167
rect -227 -1217 -223 -1167
rect -205 -1209 -201 -1169
rect -197 -1209 -193 -1169
rect -109 -1247 -105 -1167
rect -101 -1247 -97 -1167
rect -93 -1247 -89 -1167
rect -71 -1247 -67 -1167
rect -63 -1247 -59 -1167
rect -55 -1247 -51 -1167
rect -33 -1217 -29 -1167
rect -25 -1217 -21 -1167
rect 912 -1145 916 -1139
rect 921 -1145 925 -1139
rect 931 -1145 935 -1139
rect 955 -1145 959 -1139
rect 963 -1145 967 -1139
rect 711 -1167 715 -1161
rect 749 -1167 753 -1161
rect 759 -1167 763 -1161
rect 767 -1167 771 -1161
rect -3 -1209 1 -1169
rect 5 -1209 9 -1169
rect 235 -1202 239 -1196
rect 244 -1202 248 -1196
rect 254 -1202 258 -1196
rect 278 -1202 282 -1196
rect 286 -1202 290 -1196
rect 1308 -1105 1312 -1025
rect 1316 -1105 1320 -1025
rect 1324 -1105 1328 -1025
rect 1346 -1105 1350 -1025
rect 1354 -1105 1358 -1025
rect 1362 -1105 1366 -1025
rect 1384 -1075 1388 -1025
rect 1392 -1075 1396 -1025
rect 1414 -1067 1418 -1027
rect 1422 -1067 1426 -1027
rect 1509 -1067 1513 -1059
rect 1517 -1067 1521 -1059
rect 1097 -1210 1101 -1204
rect 1105 -1210 1109 -1204
rect 1113 -1210 1117 -1204
rect 1132 -1210 1136 -1204
rect 1151 -1210 1155 -1204
rect 1163 -1210 1167 -1204
rect 1171 -1210 1175 -1204
rect 526 -1221 530 -1215
rect 554 -1221 558 -1215
rect 564 -1221 568 -1215
rect 572 -1221 576 -1215
rect 911 -1236 915 -1230
rect 959 -1236 963 -1230
rect 968 -1236 972 -1230
rect 976 -1236 980 -1230
rect 235 -1277 239 -1271
rect 244 -1277 248 -1271
rect 254 -1277 258 -1271
rect 278 -1277 282 -1271
rect 286 -1277 290 -1271
rect 1309 -1294 1313 -1214
rect 1317 -1294 1321 -1214
rect 1325 -1294 1329 -1214
rect 1347 -1294 1351 -1214
rect 1355 -1294 1359 -1214
rect 1363 -1294 1367 -1214
rect 1385 -1264 1389 -1214
rect 1393 -1264 1397 -1214
rect 1415 -1256 1419 -1216
rect 1423 -1256 1427 -1216
rect 1507 -1256 1511 -1248
rect 1515 -1256 1519 -1248
rect -311 -1431 -307 -1351
rect -303 -1431 -299 -1351
rect -295 -1431 -291 -1351
rect -273 -1431 -269 -1351
rect -265 -1431 -261 -1351
rect -257 -1431 -253 -1351
rect -235 -1401 -231 -1351
rect -227 -1401 -223 -1351
rect -205 -1393 -201 -1353
rect -197 -1393 -193 -1353
rect -106 -1429 -102 -1349
rect -98 -1429 -94 -1349
rect -90 -1429 -86 -1349
rect -68 -1429 -64 -1349
rect -60 -1429 -56 -1349
rect -52 -1429 -48 -1349
rect -30 -1399 -26 -1349
rect -22 -1399 -18 -1349
rect 0 -1391 4 -1351
rect 8 -1391 12 -1351
rect 235 -1352 239 -1346
rect 244 -1352 248 -1346
rect 254 -1352 258 -1346
rect 278 -1352 282 -1346
rect 286 -1352 290 -1346
rect 1310 -1482 1314 -1402
rect 1318 -1482 1322 -1402
rect 1326 -1482 1330 -1402
rect 1348 -1482 1352 -1402
rect 1356 -1482 1360 -1402
rect 1364 -1482 1368 -1402
rect 1386 -1452 1390 -1402
rect 1394 -1452 1398 -1402
rect 1416 -1444 1420 -1404
rect 1424 -1444 1428 -1404
rect 1510 -1444 1514 -1436
rect 1518 -1444 1522 -1436
<< polysilicon >>
rect 1312 -646 1314 -636
rect 1320 -646 1322 -636
rect 1350 -646 1352 -636
rect 1358 -646 1360 -636
rect 1388 -646 1390 -636
rect 1388 -711 1390 -696
rect 1396 -711 1398 -636
rect 1418 -648 1420 -645
rect 1515 -680 1517 -677
rect 1418 -702 1420 -688
rect 231 -732 317 -730
rect 231 -740 233 -732
rect 247 -740 249 -737
rect 257 -740 259 -737
rect 267 -740 269 -732
rect 277 -740 279 -737
rect 297 -740 299 -737
rect -304 -782 -302 -772
rect -296 -782 -294 -772
rect -266 -782 -264 -772
rect -258 -782 -256 -772
rect -228 -782 -226 -772
rect -228 -847 -226 -832
rect -220 -847 -218 -772
rect -198 -784 -196 -781
rect 231 -788 233 -746
rect 247 -788 249 -746
rect 257 -767 259 -746
rect 267 -749 269 -746
rect 257 -769 269 -767
rect 257 -788 259 -785
rect 267 -788 269 -769
rect 277 -788 279 -746
rect 297 -769 299 -746
rect 315 -774 317 -732
rect 1312 -741 1314 -726
rect 1320 -733 1322 -726
rect 1350 -744 1352 -726
rect 1358 -744 1360 -726
rect 1312 -764 1314 -761
rect 288 -776 317 -774
rect -109 -802 -107 -792
rect -101 -802 -99 -792
rect -71 -802 -69 -792
rect -63 -802 -61 -792
rect -33 -802 -31 -792
rect -198 -838 -196 -824
rect -304 -877 -302 -862
rect -296 -869 -294 -862
rect -266 -880 -264 -862
rect -258 -880 -256 -862
rect -304 -900 -302 -897
rect -198 -861 -196 -858
rect -33 -867 -31 -852
rect -25 -867 -23 -792
rect 231 -795 233 -792
rect -3 -804 -1 -801
rect 247 -803 249 -792
rect 257 -798 259 -792
rect 267 -795 269 -792
rect 277 -795 279 -792
rect 288 -798 290 -776
rect 297 -788 299 -780
rect 1515 -703 1517 -688
rect 1515 -710 1517 -707
rect 1418 -725 1420 -722
rect 1388 -754 1390 -751
rect 1396 -754 1398 -751
rect 1350 -787 1352 -784
rect 1358 -787 1360 -784
rect 257 -800 290 -798
rect 297 -803 299 -792
rect 247 -805 299 -803
rect 231 -824 317 -822
rect 231 -832 233 -824
rect 247 -832 249 -829
rect 257 -832 259 -829
rect 267 -832 269 -824
rect 277 -832 279 -829
rect 297 -832 299 -829
rect -3 -858 -1 -844
rect -228 -890 -226 -887
rect -220 -890 -218 -887
rect -109 -897 -107 -882
rect -101 -889 -99 -882
rect -71 -900 -69 -882
rect -63 -900 -61 -882
rect -109 -920 -107 -917
rect -266 -923 -264 -920
rect -258 -923 -256 -920
rect -3 -881 -1 -878
rect 231 -880 233 -838
rect 247 -880 249 -838
rect 257 -859 259 -838
rect 267 -841 269 -838
rect 257 -861 269 -859
rect 257 -880 259 -877
rect 267 -880 269 -861
rect 277 -880 279 -838
rect 297 -861 299 -838
rect 315 -866 317 -824
rect 1315 -836 1317 -826
rect 1323 -836 1325 -826
rect 1353 -836 1355 -826
rect 1361 -836 1363 -826
rect 1391 -836 1393 -826
rect 919 -845 921 -836
rect 929 -845 931 -836
rect 939 -845 941 -836
rect 949 -845 951 -836
rect 959 -845 961 -836
rect 992 -845 994 -836
rect 528 -865 530 -856
rect 538 -865 540 -856
rect 571 -865 573 -856
rect 288 -868 317 -866
rect 231 -887 233 -884
rect 247 -895 249 -884
rect 257 -890 259 -884
rect 267 -887 269 -884
rect 277 -887 279 -884
rect 288 -890 290 -868
rect 297 -880 299 -872
rect 257 -892 290 -890
rect 297 -895 299 -884
rect 247 -897 299 -895
rect 528 -897 530 -871
rect 538 -897 540 -871
rect 571 -897 573 -871
rect 719 -886 721 -877
rect 729 -886 731 -877
rect 739 -886 741 -877
rect 749 -886 751 -877
rect 780 -886 782 -877
rect 528 -904 530 -901
rect 538 -904 540 -901
rect 571 -904 573 -901
rect -33 -910 -31 -907
rect -25 -910 -23 -907
rect 231 -916 317 -914
rect 231 -924 233 -916
rect 247 -924 249 -921
rect 257 -924 259 -921
rect 267 -924 269 -916
rect 277 -924 279 -921
rect 297 -924 299 -921
rect -71 -943 -69 -940
rect -63 -943 -61 -940
rect -306 -973 -304 -963
rect -298 -973 -296 -963
rect -268 -973 -266 -963
rect -260 -973 -258 -963
rect -230 -973 -228 -963
rect -230 -1038 -228 -1023
rect -222 -1038 -220 -963
rect -200 -975 -198 -972
rect 231 -972 233 -930
rect 247 -972 249 -930
rect 257 -951 259 -930
rect 267 -933 269 -930
rect 257 -953 269 -951
rect 257 -972 259 -969
rect 267 -972 269 -953
rect 277 -972 279 -930
rect 297 -953 299 -930
rect 315 -958 317 -916
rect 719 -929 721 -892
rect 729 -929 731 -892
rect 739 -929 741 -892
rect 749 -929 751 -892
rect 780 -929 782 -892
rect 919 -895 921 -851
rect 929 -895 931 -851
rect 939 -895 941 -851
rect 949 -895 951 -851
rect 959 -895 961 -851
rect 992 -895 994 -851
rect 919 -902 921 -899
rect 929 -902 931 -899
rect 939 -902 941 -899
rect 949 -902 951 -899
rect 959 -902 961 -899
rect 992 -902 994 -899
rect 1102 -900 1188 -898
rect 1102 -908 1104 -900
rect 1118 -908 1120 -905
rect 1128 -908 1130 -905
rect 1138 -908 1140 -900
rect 1148 -908 1150 -905
rect 1168 -908 1170 -905
rect 719 -936 721 -933
rect 729 -936 731 -933
rect 739 -936 741 -933
rect 749 -936 751 -933
rect 780 -936 782 -933
rect 919 -951 921 -942
rect 929 -951 931 -942
rect 939 -951 941 -942
rect 949 -951 951 -942
rect 980 -951 982 -942
rect 1102 -956 1104 -914
rect 1118 -956 1120 -914
rect 1128 -935 1130 -914
rect 1138 -917 1140 -914
rect 1128 -937 1140 -935
rect 1128 -956 1130 -953
rect 1138 -956 1140 -937
rect 1148 -956 1150 -914
rect 1168 -937 1170 -914
rect 1186 -942 1188 -900
rect 1391 -901 1393 -886
rect 1399 -901 1401 -826
rect 1421 -838 1423 -835
rect 1515 -870 1517 -867
rect 1421 -892 1423 -878
rect 1315 -931 1317 -916
rect 1323 -923 1325 -916
rect 1159 -944 1188 -942
rect 288 -960 317 -958
rect -108 -985 -106 -975
rect -100 -985 -98 -975
rect -70 -985 -68 -975
rect -62 -985 -60 -975
rect -32 -985 -30 -975
rect -200 -1029 -198 -1015
rect -306 -1068 -304 -1053
rect -298 -1060 -296 -1053
rect -268 -1071 -266 -1053
rect -260 -1071 -258 -1053
rect -306 -1091 -304 -1088
rect -200 -1052 -198 -1049
rect -32 -1050 -30 -1035
rect -24 -1050 -22 -975
rect 231 -979 233 -976
rect -2 -987 0 -984
rect 247 -987 249 -976
rect 257 -982 259 -976
rect 267 -979 269 -976
rect 277 -979 279 -976
rect 288 -982 290 -960
rect 527 -964 529 -961
rect 537 -964 539 -961
rect 555 -964 557 -961
rect 297 -972 299 -964
rect 257 -984 290 -982
rect 297 -987 299 -976
rect 247 -989 299 -987
rect 527 -1002 529 -970
rect 537 -1002 539 -970
rect 555 -1002 557 -970
rect 719 -991 721 -982
rect 729 -991 731 -982
rect 739 -991 741 -982
rect 772 -991 774 -982
rect 919 -994 921 -957
rect 929 -994 931 -957
rect 939 -994 941 -957
rect 949 -994 951 -957
rect 980 -994 982 -957
rect 1102 -963 1104 -960
rect 1118 -971 1120 -960
rect 1128 -966 1130 -960
rect 1138 -963 1140 -960
rect 1148 -963 1150 -960
rect 1159 -966 1161 -944
rect 1168 -956 1170 -948
rect 1353 -934 1355 -916
rect 1361 -934 1363 -916
rect 1315 -954 1317 -951
rect 1128 -968 1161 -966
rect 1168 -971 1170 -960
rect 1118 -973 1170 -971
rect 1515 -893 1517 -878
rect 1515 -900 1517 -897
rect 1421 -915 1423 -912
rect 1391 -944 1393 -941
rect 1399 -944 1401 -941
rect 1353 -977 1355 -974
rect 1361 -977 1363 -974
rect 231 -1009 317 -1007
rect 527 -1009 529 -1006
rect 537 -1009 539 -1006
rect 555 -1009 557 -1006
rect 231 -1017 233 -1009
rect 247 -1017 249 -1014
rect 257 -1017 259 -1014
rect 267 -1017 269 -1009
rect 277 -1017 279 -1014
rect 297 -1017 299 -1014
rect -2 -1041 0 -1027
rect -230 -1081 -228 -1078
rect -222 -1081 -220 -1078
rect -108 -1080 -106 -1065
rect -100 -1072 -98 -1065
rect -70 -1083 -68 -1065
rect -62 -1083 -60 -1065
rect -108 -1103 -106 -1100
rect -268 -1114 -266 -1111
rect -260 -1114 -258 -1111
rect -2 -1064 0 -1061
rect 231 -1065 233 -1023
rect 247 -1065 249 -1023
rect 257 -1044 259 -1023
rect 267 -1026 269 -1023
rect 257 -1046 269 -1044
rect 257 -1065 259 -1062
rect 267 -1065 269 -1046
rect 277 -1065 279 -1023
rect 297 -1046 299 -1023
rect 315 -1051 317 -1009
rect 719 -1026 721 -997
rect 729 -1026 731 -997
rect 739 -1026 741 -997
rect 772 -1026 774 -997
rect 1102 -998 1188 -996
rect 919 -1001 921 -998
rect 929 -1001 931 -998
rect 939 -1001 941 -998
rect 949 -1001 951 -998
rect 980 -1001 982 -998
rect 1102 -1006 1104 -998
rect 1118 -1006 1120 -1003
rect 1128 -1006 1130 -1003
rect 1138 -1006 1140 -998
rect 1148 -1006 1150 -1003
rect 1168 -1006 1170 -1003
rect 719 -1033 721 -1030
rect 729 -1033 731 -1030
rect 739 -1033 741 -1030
rect 772 -1033 774 -1030
rect 532 -1050 534 -1041
rect 542 -1050 544 -1041
rect 552 -1050 554 -1041
rect 585 -1050 587 -1041
rect 288 -1053 317 -1051
rect 231 -1072 233 -1069
rect 247 -1080 249 -1069
rect 257 -1075 259 -1069
rect 267 -1072 269 -1069
rect 277 -1072 279 -1069
rect 288 -1075 290 -1053
rect 919 -1052 921 -1043
rect 929 -1052 931 -1043
rect 939 -1052 941 -1043
rect 972 -1052 974 -1043
rect 297 -1065 299 -1057
rect 257 -1077 290 -1075
rect 297 -1080 299 -1069
rect 247 -1082 299 -1080
rect 532 -1085 534 -1056
rect 542 -1085 544 -1056
rect 552 -1085 554 -1056
rect 585 -1085 587 -1056
rect 1102 -1054 1104 -1012
rect 1118 -1054 1120 -1012
rect 1128 -1033 1130 -1012
rect 1138 -1015 1140 -1012
rect 1128 -1035 1140 -1033
rect 1128 -1054 1130 -1051
rect 1138 -1054 1140 -1035
rect 1148 -1054 1150 -1012
rect 1168 -1035 1170 -1012
rect 1186 -1040 1188 -998
rect 1313 -1025 1315 -1015
rect 1321 -1025 1323 -1015
rect 1351 -1025 1353 -1015
rect 1359 -1025 1361 -1015
rect 1389 -1025 1391 -1015
rect 1159 -1042 1188 -1040
rect 718 -1082 720 -1073
rect 728 -1082 730 -1073
rect 761 -1082 763 -1073
rect 919 -1087 921 -1058
rect 929 -1087 931 -1058
rect 939 -1087 941 -1058
rect 972 -1087 974 -1058
rect 1102 -1061 1104 -1058
rect 1118 -1069 1120 -1058
rect 1128 -1064 1130 -1058
rect 1138 -1061 1140 -1058
rect 1148 -1061 1150 -1058
rect 1159 -1064 1161 -1042
rect 1168 -1054 1170 -1046
rect 1128 -1066 1161 -1064
rect 1168 -1069 1170 -1058
rect 1118 -1071 1170 -1069
rect -32 -1093 -30 -1090
rect -24 -1093 -22 -1090
rect 532 -1092 534 -1089
rect 542 -1092 544 -1089
rect 552 -1092 554 -1089
rect 585 -1092 587 -1089
rect 241 -1121 243 -1112
rect 251 -1121 253 -1112
rect 284 -1121 286 -1112
rect 718 -1114 720 -1088
rect 728 -1114 730 -1088
rect 761 -1114 763 -1088
rect 919 -1094 921 -1091
rect 929 -1094 931 -1091
rect 939 -1094 941 -1091
rect 972 -1094 974 -1091
rect 1102 -1098 1188 -1096
rect 1102 -1106 1104 -1098
rect 1118 -1106 1120 -1103
rect 1128 -1106 1130 -1103
rect 1138 -1106 1140 -1098
rect 1148 -1106 1150 -1103
rect 1168 -1106 1170 -1103
rect 718 -1121 720 -1118
rect 728 -1121 730 -1118
rect 761 -1121 763 -1118
rect -70 -1126 -68 -1123
rect -62 -1126 -60 -1123
rect 241 -1153 243 -1127
rect 251 -1153 253 -1127
rect 284 -1153 286 -1127
rect 532 -1136 534 -1127
rect 542 -1136 544 -1127
rect 575 -1136 577 -1127
rect 917 -1139 919 -1130
rect 927 -1139 929 -1130
rect 960 -1139 962 -1130
rect -306 -1167 -304 -1157
rect -298 -1167 -296 -1157
rect -268 -1167 -266 -1157
rect -260 -1167 -258 -1157
rect -230 -1167 -228 -1157
rect -230 -1232 -228 -1217
rect -222 -1232 -220 -1157
rect -200 -1169 -198 -1166
rect -104 -1167 -102 -1157
rect -96 -1167 -94 -1157
rect -66 -1167 -64 -1157
rect -58 -1167 -56 -1157
rect -28 -1167 -26 -1157
rect -200 -1223 -198 -1209
rect -306 -1262 -304 -1247
rect -298 -1254 -296 -1247
rect -268 -1265 -266 -1247
rect -260 -1265 -258 -1247
rect -306 -1285 -304 -1282
rect -200 -1246 -198 -1243
rect -28 -1232 -26 -1217
rect -20 -1232 -18 -1157
rect 241 -1160 243 -1157
rect 251 -1160 253 -1157
rect 284 -1160 286 -1157
rect 2 -1169 4 -1166
rect 532 -1168 534 -1142
rect 542 -1168 544 -1142
rect 575 -1168 577 -1142
rect 716 -1161 718 -1158
rect 726 -1161 728 -1158
rect 735 -1161 737 -1158
rect 745 -1161 747 -1158
rect 764 -1161 766 -1158
rect 532 -1175 534 -1172
rect 542 -1175 544 -1172
rect 575 -1175 577 -1172
rect 240 -1196 242 -1187
rect 250 -1196 252 -1187
rect 283 -1196 285 -1187
rect 2 -1223 4 -1209
rect -104 -1262 -102 -1247
rect -96 -1254 -94 -1247
rect -230 -1275 -228 -1272
rect -222 -1275 -220 -1272
rect -66 -1265 -64 -1247
rect -58 -1265 -56 -1247
rect -104 -1285 -102 -1282
rect 240 -1228 242 -1202
rect 250 -1228 252 -1202
rect 283 -1228 285 -1202
rect 531 -1215 533 -1212
rect 541 -1215 543 -1212
rect 550 -1215 552 -1212
rect 569 -1215 571 -1212
rect 716 -1213 718 -1167
rect 726 -1213 728 -1167
rect 735 -1190 737 -1167
rect 736 -1194 737 -1190
rect 735 -1213 737 -1194
rect 745 -1213 747 -1167
rect 764 -1213 766 -1167
rect 917 -1171 919 -1145
rect 927 -1171 929 -1145
rect 960 -1171 962 -1145
rect 1102 -1154 1104 -1112
rect 1118 -1154 1120 -1112
rect 1128 -1133 1130 -1112
rect 1138 -1115 1140 -1112
rect 1128 -1135 1140 -1133
rect 1128 -1154 1130 -1151
rect 1138 -1154 1140 -1135
rect 1148 -1154 1150 -1112
rect 1168 -1135 1170 -1112
rect 1186 -1140 1188 -1098
rect 1389 -1090 1391 -1075
rect 1397 -1090 1399 -1015
rect 1419 -1027 1421 -1024
rect 1514 -1059 1516 -1056
rect 1419 -1081 1421 -1067
rect 1313 -1120 1315 -1105
rect 1321 -1112 1323 -1105
rect 1351 -1123 1353 -1105
rect 1359 -1123 1361 -1105
rect 1159 -1142 1188 -1140
rect 1102 -1161 1104 -1158
rect 1118 -1169 1120 -1158
rect 1128 -1164 1130 -1158
rect 1138 -1161 1140 -1158
rect 1148 -1161 1150 -1158
rect 1159 -1164 1161 -1142
rect 1313 -1143 1315 -1140
rect 1168 -1154 1170 -1146
rect 1128 -1166 1161 -1164
rect 1168 -1169 1170 -1158
rect 1514 -1082 1516 -1067
rect 1514 -1089 1516 -1086
rect 1419 -1104 1421 -1101
rect 1389 -1133 1391 -1130
rect 1397 -1133 1399 -1130
rect 1351 -1166 1353 -1163
rect 1359 -1166 1361 -1163
rect 1118 -1171 1170 -1169
rect 917 -1178 919 -1175
rect 927 -1178 929 -1175
rect 960 -1178 962 -1175
rect 1102 -1196 1188 -1194
rect 1102 -1204 1104 -1196
rect 1118 -1204 1120 -1201
rect 1128 -1204 1130 -1201
rect 1138 -1204 1140 -1196
rect 1148 -1204 1150 -1201
rect 1168 -1204 1170 -1201
rect 716 -1220 718 -1217
rect 726 -1220 728 -1217
rect 735 -1220 737 -1217
rect 745 -1220 747 -1217
rect 764 -1220 766 -1217
rect 240 -1235 242 -1232
rect 250 -1235 252 -1232
rect 283 -1235 285 -1232
rect 2 -1246 4 -1243
rect 531 -1260 533 -1221
rect 541 -1260 543 -1221
rect 550 -1244 552 -1221
rect 551 -1248 552 -1244
rect 550 -1260 552 -1248
rect 569 -1260 571 -1221
rect 916 -1230 918 -1227
rect 926 -1230 928 -1227
rect 935 -1230 937 -1227
rect 945 -1230 947 -1227
rect 955 -1230 957 -1227
rect 973 -1230 975 -1227
rect 240 -1271 242 -1262
rect 250 -1271 252 -1262
rect 283 -1271 285 -1262
rect 531 -1267 533 -1264
rect 541 -1267 543 -1264
rect 550 -1267 552 -1264
rect 569 -1267 571 -1264
rect -28 -1275 -26 -1272
rect -20 -1275 -18 -1272
rect 240 -1303 242 -1277
rect 250 -1303 252 -1277
rect 283 -1303 285 -1277
rect 916 -1289 918 -1236
rect 926 -1289 928 -1236
rect 935 -1259 937 -1236
rect 936 -1263 937 -1259
rect 935 -1289 937 -1263
rect 945 -1289 947 -1236
rect 955 -1289 957 -1236
rect 973 -1289 975 -1236
rect 1102 -1252 1104 -1210
rect 1118 -1252 1120 -1210
rect 1128 -1231 1130 -1210
rect 1138 -1213 1140 -1210
rect 1128 -1233 1140 -1231
rect 1128 -1252 1130 -1249
rect 1138 -1252 1140 -1233
rect 1148 -1252 1150 -1210
rect 1168 -1233 1170 -1210
rect 1186 -1238 1188 -1196
rect 1314 -1214 1316 -1204
rect 1322 -1214 1324 -1204
rect 1352 -1214 1354 -1204
rect 1360 -1214 1362 -1204
rect 1390 -1214 1392 -1204
rect 1159 -1240 1188 -1238
rect 1102 -1259 1104 -1256
rect 1118 -1267 1120 -1256
rect 1128 -1262 1130 -1256
rect 1138 -1259 1140 -1256
rect 1148 -1259 1150 -1256
rect 1159 -1262 1161 -1240
rect 1168 -1252 1170 -1244
rect 1128 -1264 1161 -1262
rect 1168 -1267 1170 -1256
rect 1118 -1269 1170 -1267
rect 916 -1296 918 -1293
rect 926 -1296 928 -1293
rect 935 -1296 937 -1293
rect 945 -1296 947 -1293
rect 955 -1296 957 -1293
rect 973 -1296 975 -1293
rect 1390 -1279 1392 -1264
rect 1398 -1279 1400 -1204
rect 1420 -1216 1422 -1213
rect 1512 -1248 1514 -1245
rect 1420 -1270 1422 -1256
rect -268 -1308 -266 -1305
rect -260 -1308 -258 -1305
rect -66 -1308 -64 -1305
rect -58 -1308 -56 -1305
rect 240 -1310 242 -1307
rect 250 -1310 252 -1307
rect 283 -1310 285 -1307
rect 1314 -1309 1316 -1294
rect 1322 -1301 1324 -1294
rect 1352 -1312 1354 -1294
rect 1360 -1312 1362 -1294
rect 1314 -1332 1316 -1329
rect -306 -1351 -304 -1341
rect -298 -1351 -296 -1341
rect -268 -1351 -266 -1341
rect -260 -1351 -258 -1341
rect -230 -1351 -228 -1341
rect -230 -1416 -228 -1401
rect -222 -1416 -220 -1341
rect -101 -1349 -99 -1339
rect -93 -1349 -91 -1339
rect -63 -1349 -61 -1339
rect -55 -1349 -53 -1339
rect -25 -1349 -23 -1339
rect -200 -1353 -198 -1350
rect -200 -1407 -198 -1393
rect -306 -1446 -304 -1431
rect -298 -1438 -296 -1431
rect -268 -1449 -266 -1431
rect -260 -1449 -258 -1431
rect -306 -1469 -304 -1466
rect -200 -1430 -198 -1427
rect -25 -1414 -23 -1399
rect -17 -1414 -15 -1339
rect 240 -1346 242 -1337
rect 250 -1346 252 -1337
rect 283 -1346 285 -1337
rect 5 -1351 7 -1348
rect 1512 -1271 1514 -1256
rect 1512 -1278 1514 -1275
rect 1420 -1293 1422 -1290
rect 1390 -1322 1392 -1319
rect 1398 -1322 1400 -1319
rect 240 -1378 242 -1352
rect 250 -1378 252 -1352
rect 283 -1378 285 -1352
rect 1352 -1355 1354 -1352
rect 1360 -1355 1362 -1352
rect 240 -1385 242 -1382
rect 250 -1385 252 -1382
rect 283 -1385 285 -1382
rect 5 -1405 7 -1391
rect 1315 -1402 1317 -1392
rect 1323 -1402 1325 -1392
rect 1353 -1402 1355 -1392
rect 1361 -1402 1363 -1392
rect 1391 -1402 1393 -1392
rect -101 -1444 -99 -1429
rect -93 -1436 -91 -1429
rect -230 -1459 -228 -1456
rect -222 -1459 -220 -1456
rect -63 -1447 -61 -1429
rect -55 -1447 -53 -1429
rect -101 -1467 -99 -1464
rect 5 -1428 7 -1425
rect -25 -1457 -23 -1454
rect -17 -1457 -15 -1454
rect 1391 -1467 1393 -1452
rect 1399 -1467 1401 -1392
rect 1421 -1404 1423 -1401
rect 1515 -1436 1517 -1433
rect 1421 -1458 1423 -1444
rect -268 -1492 -266 -1489
rect -260 -1492 -258 -1489
rect -63 -1490 -61 -1487
rect -55 -1490 -53 -1487
rect 1315 -1497 1317 -1482
rect 1323 -1489 1325 -1482
rect 1353 -1500 1355 -1482
rect 1361 -1500 1363 -1482
rect 1315 -1520 1317 -1517
rect 1515 -1459 1517 -1444
rect 1515 -1466 1517 -1463
rect 1421 -1481 1423 -1478
rect 1391 -1510 1393 -1507
rect 1399 -1510 1401 -1507
rect 1353 -1543 1355 -1540
rect 1361 -1543 1363 -1540
<< polycontact >>
rect 1311 -636 1315 -632
rect 1319 -636 1323 -632
rect 1349 -636 1353 -632
rect 1357 -636 1361 -632
rect 1387 -636 1391 -632
rect 1395 -636 1399 -632
rect 1414 -699 1418 -695
rect 1511 -700 1515 -696
rect -305 -772 -301 -768
rect -297 -772 -293 -768
rect -267 -772 -263 -768
rect -259 -772 -255 -768
rect -229 -772 -225 -768
rect -221 -772 -217 -768
rect 227 -769 231 -765
rect 253 -769 257 -765
rect 279 -769 283 -765
rect 299 -769 303 -765
rect -110 -792 -106 -788
rect -102 -792 -98 -788
rect -72 -792 -68 -788
rect -64 -792 -60 -788
rect -34 -792 -30 -788
rect -26 -792 -22 -788
rect -202 -835 -198 -831
rect 299 -784 303 -780
rect -7 -855 -3 -851
rect 227 -861 231 -857
rect 253 -861 257 -857
rect 279 -861 283 -857
rect 299 -861 303 -857
rect 1314 -826 1318 -822
rect 1322 -826 1326 -822
rect 1352 -826 1356 -822
rect 1360 -826 1364 -822
rect 1390 -826 1394 -822
rect 1398 -826 1402 -822
rect 915 -863 919 -859
rect 299 -876 303 -872
rect 524 -883 528 -879
rect 534 -892 538 -888
rect 567 -883 571 -879
rect 715 -904 719 -900
rect 227 -953 231 -949
rect -307 -963 -303 -959
rect -299 -963 -295 -959
rect -269 -963 -265 -959
rect -261 -963 -257 -959
rect -231 -963 -227 -959
rect -223 -963 -219 -959
rect -109 -975 -105 -971
rect -101 -975 -97 -971
rect -71 -975 -67 -971
rect -63 -975 -59 -971
rect -33 -975 -29 -971
rect -25 -975 -21 -971
rect 253 -953 257 -949
rect 279 -953 283 -949
rect 299 -953 303 -949
rect 725 -911 729 -907
rect 735 -918 739 -914
rect 745 -925 749 -921
rect 776 -904 780 -900
rect 925 -870 929 -866
rect 935 -877 939 -873
rect 945 -884 949 -880
rect 955 -892 959 -888
rect 988 -863 992 -859
rect 1098 -937 1102 -933
rect 1124 -937 1128 -933
rect 1150 -937 1154 -933
rect 1170 -937 1174 -933
rect 1417 -889 1421 -885
rect 1511 -890 1515 -886
rect -204 -1026 -200 -1022
rect 299 -968 303 -964
rect 915 -969 919 -965
rect 523 -983 527 -979
rect 533 -990 537 -986
rect 551 -988 555 -984
rect 925 -976 929 -972
rect 935 -983 939 -979
rect 945 -990 949 -986
rect 976 -969 980 -965
rect 1170 -952 1174 -948
rect 715 -1009 719 -1005
rect -6 -1038 -2 -1034
rect 227 -1046 231 -1042
rect 253 -1046 257 -1042
rect 279 -1046 283 -1042
rect 299 -1046 303 -1042
rect 725 -1016 729 -1012
rect 735 -1023 739 -1019
rect 768 -1009 772 -1005
rect 1098 -1035 1102 -1031
rect 299 -1061 303 -1057
rect 528 -1068 532 -1064
rect 538 -1075 542 -1071
rect 548 -1082 552 -1078
rect 581 -1068 585 -1064
rect 1124 -1035 1128 -1031
rect 1150 -1035 1154 -1031
rect 1170 -1035 1174 -1031
rect 1312 -1015 1316 -1011
rect 1320 -1015 1324 -1011
rect 1350 -1015 1354 -1011
rect 1358 -1015 1362 -1011
rect 1388 -1015 1392 -1011
rect 1396 -1015 1400 -1011
rect 915 -1070 919 -1066
rect 925 -1077 929 -1073
rect 935 -1084 939 -1080
rect 968 -1070 972 -1066
rect 1170 -1050 1174 -1046
rect 714 -1100 718 -1096
rect 724 -1109 728 -1105
rect 757 -1100 761 -1096
rect 237 -1139 241 -1135
rect 247 -1148 251 -1144
rect 280 -1139 284 -1135
rect 1098 -1135 1102 -1131
rect -307 -1157 -303 -1153
rect -299 -1157 -295 -1153
rect -269 -1157 -265 -1153
rect -261 -1157 -257 -1153
rect -231 -1157 -227 -1153
rect -223 -1157 -219 -1153
rect -105 -1157 -101 -1153
rect -97 -1157 -93 -1153
rect -67 -1157 -63 -1153
rect -59 -1157 -55 -1153
rect -29 -1157 -25 -1153
rect -21 -1157 -17 -1153
rect 528 -1154 532 -1150
rect -204 -1220 -200 -1216
rect 538 -1163 542 -1159
rect 571 -1154 575 -1150
rect 913 -1157 917 -1153
rect 712 -1180 716 -1176
rect -2 -1220 2 -1216
rect 236 -1214 240 -1210
rect 246 -1223 250 -1219
rect 279 -1214 283 -1210
rect 722 -1187 726 -1183
rect 732 -1194 736 -1190
rect 741 -1201 745 -1197
rect 760 -1185 764 -1181
rect 923 -1166 927 -1162
rect 956 -1157 960 -1153
rect 1124 -1135 1128 -1131
rect 1150 -1135 1154 -1131
rect 1170 -1135 1174 -1131
rect 1415 -1078 1419 -1074
rect 1510 -1079 1514 -1075
rect 1170 -1150 1174 -1146
rect 527 -1234 531 -1230
rect 537 -1241 541 -1237
rect 565 -1239 569 -1235
rect 547 -1248 551 -1244
rect 1098 -1233 1102 -1229
rect 912 -1249 916 -1245
rect 236 -1289 240 -1285
rect 246 -1298 250 -1294
rect 279 -1289 283 -1285
rect 922 -1256 926 -1252
rect 932 -1263 936 -1259
rect 941 -1270 945 -1266
rect 951 -1277 955 -1273
rect 969 -1254 973 -1250
rect 1124 -1233 1128 -1229
rect 1150 -1233 1154 -1229
rect 1170 -1233 1174 -1229
rect 1313 -1204 1317 -1200
rect 1321 -1204 1325 -1200
rect 1351 -1204 1355 -1200
rect 1359 -1204 1363 -1200
rect 1389 -1204 1393 -1200
rect 1397 -1204 1401 -1200
rect 1170 -1248 1174 -1244
rect 1416 -1267 1420 -1263
rect 1508 -1268 1512 -1264
rect -307 -1341 -303 -1337
rect -299 -1341 -295 -1337
rect -269 -1341 -265 -1337
rect -261 -1341 -257 -1337
rect -231 -1341 -227 -1337
rect -223 -1341 -219 -1337
rect -102 -1339 -98 -1335
rect -94 -1339 -90 -1335
rect -64 -1339 -60 -1335
rect -56 -1339 -52 -1335
rect -26 -1339 -22 -1335
rect -18 -1339 -14 -1335
rect -204 -1404 -200 -1400
rect 236 -1364 240 -1360
rect 246 -1373 250 -1369
rect 279 -1364 283 -1360
rect 1 -1402 5 -1398
rect 1314 -1392 1318 -1388
rect 1322 -1392 1326 -1388
rect 1352 -1392 1356 -1388
rect 1360 -1392 1364 -1388
rect 1390 -1392 1394 -1388
rect 1398 -1392 1402 -1388
rect 1417 -1455 1421 -1451
rect 1511 -1456 1515 -1452
<< metal1 >>
rect -381 -535 1500 -502
rect -297 -757 -278 -535
rect 1319 -625 1399 -621
rect 1311 -632 1315 -628
rect 1319 -632 1323 -625
rect 1335 -632 1353 -628
rect 1310 -645 1311 -639
rect 1307 -646 1311 -645
rect 218 -727 419 -723
rect 218 -731 230 -727
rect 226 -740 230 -731
rect 242 -740 246 -727
rect 280 -740 284 -727
rect 300 -728 419 -727
rect 300 -740 304 -728
rect -297 -761 -217 -757
rect -305 -768 -301 -764
rect -297 -768 -293 -761
rect -281 -768 -263 -764
rect -306 -781 -305 -775
rect -309 -782 -305 -781
rect -293 -871 -289 -862
rect -281 -871 -277 -768
rect -259 -768 -255 -761
rect -245 -768 -225 -764
rect -255 -781 -253 -777
rect -255 -782 -250 -781
rect -309 -874 -277 -871
rect -271 -872 -267 -862
rect -245 -872 -241 -768
rect -221 -768 -217 -761
rect -183 -765 179 -762
rect 234 -765 238 -746
rect 261 -756 265 -746
rect -183 -769 227 -765
rect 234 -769 253 -765
rect -233 -780 -229 -777
rect -206 -780 -185 -775
rect -238 -781 -229 -780
rect -233 -782 -229 -781
rect -203 -784 -199 -780
rect -221 -831 -213 -829
rect -221 -832 -202 -831
rect -217 -835 -202 -832
rect -195 -832 -191 -824
rect -182 -832 -176 -769
rect 15 -777 220 -772
rect 225 -777 227 -773
rect -102 -781 -22 -777
rect -110 -788 -106 -784
rect -102 -788 -98 -781
rect -86 -788 -68 -784
rect -111 -801 -110 -795
rect -217 -847 -213 -835
rect -195 -836 -176 -832
rect -114 -802 -110 -801
rect -195 -838 -191 -836
rect -309 -877 -305 -874
rect -271 -877 -241 -872
rect -301 -929 -297 -897
rect -271 -880 -267 -877
rect -255 -922 -251 -920
rect -203 -867 -199 -858
rect -209 -871 -185 -867
rect -233 -893 -229 -887
rect -209 -893 -206 -871
rect -98 -891 -94 -882
rect -86 -891 -82 -788
rect -64 -788 -60 -781
rect -50 -788 -30 -784
rect -60 -801 -58 -797
rect -60 -802 -55 -801
rect -233 -897 -206 -893
rect -114 -894 -82 -891
rect -76 -892 -72 -882
rect -50 -892 -46 -788
rect -26 -788 -22 -781
rect -38 -800 -34 -797
rect -11 -800 10 -795
rect -43 -801 -34 -800
rect -38 -802 -34 -801
rect -8 -804 -4 -800
rect -26 -851 -18 -849
rect -26 -852 -7 -851
rect -22 -855 -7 -852
rect 0 -852 4 -844
rect 15 -852 19 -777
rect 112 -779 119 -777
rect 234 -788 238 -769
rect 261 -788 265 -761
rect 292 -765 296 -746
rect 336 -756 343 -741
rect 327 -761 343 -756
rect 283 -769 296 -765
rect 292 -788 296 -769
rect 303 -772 307 -765
rect 303 -784 307 -777
rect 226 -806 230 -792
rect 242 -806 246 -792
rect 280 -806 284 -792
rect 300 -806 304 -792
rect 226 -810 311 -806
rect 218 -819 310 -815
rect 218 -823 230 -819
rect 226 -832 230 -823
rect 242 -832 246 -819
rect 280 -832 284 -819
rect 300 -832 304 -819
rect -22 -867 -18 -855
rect 0 -856 19 -852
rect 0 -858 4 -856
rect -114 -897 -110 -894
rect -76 -897 -46 -892
rect -233 -922 -229 -897
rect -255 -926 -229 -922
rect -255 -929 -251 -926
rect -301 -933 -251 -929
rect -299 -952 -219 -948
rect -307 -959 -303 -955
rect -299 -959 -295 -952
rect -283 -959 -265 -955
rect -308 -972 -307 -966
rect -311 -973 -307 -972
rect -295 -1062 -291 -1053
rect -283 -1062 -279 -959
rect -261 -959 -257 -952
rect -247 -959 -227 -955
rect -257 -972 -255 -968
rect -257 -973 -252 -972
rect -311 -1065 -279 -1062
rect -273 -1063 -269 -1053
rect -247 -1063 -243 -959
rect -223 -959 -219 -952
rect -106 -949 -102 -917
rect -76 -900 -72 -897
rect -60 -942 -56 -940
rect 24 -857 166 -854
rect 234 -857 238 -838
rect 261 -848 265 -838
rect 24 -861 227 -857
rect 234 -861 253 -857
rect 24 -862 31 -861
rect 53 -865 220 -864
rect 24 -869 220 -865
rect -8 -887 -4 -878
rect -14 -891 10 -887
rect -38 -913 -34 -907
rect -14 -913 -11 -891
rect -38 -917 -11 -913
rect -38 -942 -34 -917
rect -60 -946 -34 -942
rect -60 -949 -56 -946
rect -106 -953 -56 -949
rect -101 -964 -21 -960
rect -235 -971 -231 -968
rect -208 -971 -187 -966
rect -109 -971 -105 -967
rect -240 -972 -231 -971
rect -235 -973 -231 -972
rect -205 -975 -201 -971
rect -101 -971 -97 -964
rect -85 -971 -67 -967
rect -110 -984 -109 -978
rect -223 -1022 -215 -1020
rect -223 -1023 -204 -1022
rect -219 -1026 -204 -1023
rect -197 -1023 -193 -1015
rect -113 -985 -109 -984
rect -219 -1038 -215 -1026
rect -197 -1027 -180 -1023
rect -197 -1029 -193 -1027
rect -311 -1068 -307 -1065
rect -273 -1068 -243 -1063
rect -303 -1120 -299 -1088
rect -273 -1071 -269 -1068
rect -257 -1113 -253 -1111
rect -205 -1058 -201 -1049
rect -211 -1062 -187 -1058
rect -235 -1084 -231 -1078
rect -211 -1084 -208 -1062
rect -97 -1074 -93 -1065
rect -85 -1074 -81 -971
rect -63 -971 -59 -964
rect -49 -971 -29 -967
rect -59 -984 -57 -980
rect -59 -985 -54 -984
rect -235 -1088 -208 -1084
rect -113 -1077 -81 -1074
rect -75 -1075 -71 -1065
rect -49 -1075 -45 -971
rect -25 -971 -21 -964
rect -37 -983 -33 -980
rect -10 -983 11 -978
rect -42 -984 -33 -983
rect -37 -985 -33 -984
rect -7 -987 -3 -983
rect -25 -1034 -17 -1032
rect -25 -1035 -6 -1034
rect -21 -1038 -6 -1035
rect 1 -1035 5 -1027
rect 24 -1035 31 -869
rect 101 -871 108 -869
rect 234 -880 238 -861
rect 261 -880 265 -853
rect 292 -857 296 -838
rect 358 -848 364 -779
rect 327 -853 364 -848
rect 413 -846 419 -728
rect 1323 -735 1327 -726
rect 1335 -735 1339 -632
rect 1357 -632 1361 -625
rect 1371 -632 1391 -628
rect 1361 -645 1363 -641
rect 1361 -646 1366 -645
rect 1307 -738 1339 -735
rect 1345 -736 1349 -726
rect 1371 -736 1375 -632
rect 1395 -632 1399 -625
rect 1383 -644 1387 -641
rect 1410 -644 1510 -639
rect 1378 -645 1387 -644
rect 1383 -646 1387 -645
rect 1413 -648 1417 -644
rect 1503 -672 1510 -644
rect 1503 -676 1528 -672
rect 1510 -680 1514 -676
rect 1395 -695 1403 -693
rect 1395 -696 1414 -695
rect 1399 -699 1414 -696
rect 1421 -696 1425 -688
rect 1518 -696 1522 -688
rect 1399 -711 1403 -699
rect 1421 -700 1511 -696
rect 1518 -700 1531 -696
rect 1421 -702 1425 -700
rect 1307 -741 1311 -738
rect 1345 -741 1375 -736
rect 1315 -793 1319 -761
rect 1345 -744 1349 -741
rect 1361 -786 1365 -784
rect 1518 -703 1522 -700
rect 1510 -711 1514 -707
rect 1503 -715 1528 -711
rect 1413 -731 1417 -722
rect 1503 -730 1509 -715
rect 1431 -731 1509 -730
rect 1407 -735 1509 -731
rect 1383 -757 1387 -751
rect 1407 -757 1410 -735
rect 1383 -761 1410 -757
rect 1383 -786 1387 -761
rect 1361 -790 1387 -786
rect 1361 -793 1365 -790
rect 1315 -797 1365 -793
rect 1322 -815 1402 -811
rect 619 -828 882 -821
rect 1314 -822 1318 -818
rect 1322 -822 1326 -815
rect 1338 -822 1356 -818
rect 578 -846 586 -845
rect 413 -850 586 -846
rect 413 -851 528 -850
rect 283 -861 296 -857
rect 292 -880 296 -861
rect 303 -864 307 -857
rect 303 -876 307 -869
rect 523 -865 527 -851
rect 542 -865 546 -850
rect 566 -865 570 -850
rect 578 -853 586 -850
rect 877 -866 882 -828
rect 907 -830 1004 -826
rect 907 -834 918 -830
rect 914 -845 918 -834
rect 933 -845 937 -830
rect 953 -845 957 -830
rect 987 -845 991 -830
rect 1313 -835 1314 -829
rect 1310 -836 1314 -835
rect 897 -859 913 -858
rect 923 -859 927 -851
rect 943 -859 947 -851
rect 963 -859 967 -851
rect 995 -859 999 -851
rect 897 -863 915 -859
rect 923 -863 988 -859
rect 995 -863 1016 -859
rect 386 -883 471 -879
rect 532 -879 536 -871
rect 574 -879 578 -871
rect 706 -871 793 -867
rect 877 -870 925 -866
rect 706 -875 718 -871
rect 482 -882 524 -879
rect 475 -883 524 -882
rect 532 -883 567 -879
rect 574 -883 603 -879
rect 386 -884 391 -883
rect 444 -884 450 -883
rect 226 -894 230 -884
rect 222 -898 230 -894
rect 242 -898 246 -884
rect 280 -898 284 -884
rect 300 -898 304 -884
rect 464 -885 471 -883
rect 400 -892 534 -888
rect 400 -893 405 -892
rect 542 -897 546 -883
rect 574 -897 578 -883
rect 594 -884 603 -883
rect 714 -886 718 -875
rect 733 -886 737 -871
rect 753 -886 757 -871
rect 775 -886 779 -871
rect 853 -877 935 -873
rect 817 -884 945 -880
rect 817 -885 920 -884
rect 817 -886 824 -885
rect 222 -902 311 -898
rect 218 -911 310 -907
rect 523 -908 527 -901
rect 566 -908 570 -901
rect 723 -900 727 -892
rect 743 -900 747 -892
rect 783 -900 787 -892
rect 835 -892 955 -888
rect 835 -893 841 -892
rect 963 -895 967 -863
rect 995 -895 999 -863
rect 1011 -864 1016 -863
rect 1098 -895 1181 -891
rect 642 -904 715 -900
rect 723 -904 776 -900
rect 783 -904 806 -900
rect 218 -915 230 -911
rect 226 -924 230 -915
rect 242 -924 246 -911
rect 280 -924 284 -911
rect 300 -924 304 -911
rect 516 -912 585 -908
rect 620 -911 725 -907
rect 620 -918 735 -914
rect 620 -920 626 -918
rect 632 -925 745 -921
rect 632 -926 639 -925
rect 753 -929 757 -904
rect 783 -929 787 -904
rect 801 -905 806 -904
rect 914 -906 918 -899
rect 987 -906 991 -899
rect 1098 -900 1101 -895
rect 1001 -906 1009 -903
rect 907 -910 1009 -906
rect 1097 -908 1101 -900
rect 1113 -908 1117 -895
rect 1151 -908 1155 -895
rect 1171 -908 1175 -895
rect 53 -949 153 -946
rect 234 -949 238 -930
rect 261 -940 265 -930
rect 53 -953 227 -949
rect 234 -953 253 -949
rect -21 -1050 -17 -1038
rect 1 -1039 31 -1035
rect 35 -961 220 -956
rect 1 -1041 5 -1039
rect -113 -1080 -109 -1077
rect -75 -1080 -45 -1075
rect -235 -1113 -231 -1088
rect -257 -1117 -231 -1113
rect -257 -1120 -253 -1117
rect -303 -1124 -253 -1120
rect -105 -1129 -101 -1100
rect -75 -1083 -71 -1080
rect -106 -1132 -101 -1129
rect -59 -1125 -55 -1123
rect -7 -1070 -3 -1061
rect -13 -1074 11 -1070
rect -37 -1096 -33 -1090
rect -13 -1096 -10 -1074
rect -37 -1100 -10 -1096
rect -37 -1125 -33 -1100
rect -59 -1129 -33 -1125
rect -59 -1132 -55 -1129
rect -106 -1136 -55 -1132
rect -106 -1138 -102 -1136
rect -299 -1146 -219 -1142
rect -307 -1153 -303 -1149
rect -299 -1153 -295 -1146
rect -283 -1153 -265 -1149
rect -308 -1166 -307 -1160
rect -311 -1167 -307 -1166
rect -295 -1256 -291 -1247
rect -283 -1256 -279 -1153
rect -261 -1153 -257 -1146
rect -247 -1153 -227 -1149
rect -257 -1166 -255 -1162
rect -257 -1167 -252 -1166
rect -311 -1259 -279 -1256
rect -273 -1257 -269 -1247
rect -247 -1257 -243 -1153
rect -223 -1153 -219 -1146
rect -97 -1146 -17 -1142
rect -105 -1153 -101 -1149
rect -97 -1153 -93 -1146
rect -81 -1153 -63 -1149
rect -235 -1165 -231 -1162
rect -208 -1165 -187 -1160
rect -240 -1166 -231 -1165
rect -235 -1167 -231 -1166
rect -205 -1169 -201 -1165
rect -106 -1166 -105 -1160
rect -109 -1167 -105 -1166
rect -223 -1216 -215 -1214
rect -223 -1217 -204 -1216
rect -219 -1220 -204 -1217
rect -197 -1217 -193 -1209
rect -219 -1232 -215 -1220
rect -197 -1221 -178 -1217
rect -197 -1223 -193 -1221
rect -311 -1262 -307 -1259
rect -273 -1262 -243 -1257
rect -303 -1314 -299 -1282
rect -273 -1265 -269 -1262
rect -257 -1307 -253 -1305
rect -205 -1252 -201 -1243
rect -211 -1256 -187 -1252
rect -93 -1256 -89 -1247
rect -81 -1256 -77 -1153
rect -59 -1153 -55 -1146
rect -45 -1153 -25 -1149
rect -55 -1166 -53 -1162
rect -55 -1167 -50 -1166
rect -235 -1278 -231 -1272
rect -211 -1278 -208 -1256
rect -235 -1282 -208 -1278
rect -109 -1259 -77 -1256
rect -71 -1257 -67 -1247
rect -45 -1257 -41 -1153
rect -21 -1153 -17 -1146
rect -33 -1165 -29 -1162
rect -6 -1165 15 -1160
rect -38 -1166 -29 -1165
rect -33 -1167 -29 -1166
rect -3 -1169 1 -1165
rect -21 -1216 -13 -1214
rect -21 -1217 -2 -1216
rect -17 -1220 -2 -1217
rect 5 -1217 9 -1209
rect 35 -1217 39 -961
rect 89 -963 96 -961
rect 234 -972 238 -953
rect 261 -972 265 -945
rect 292 -949 296 -930
rect 327 -945 378 -940
rect 464 -942 592 -935
rect 714 -938 718 -933
rect 283 -953 296 -949
rect 292 -972 296 -953
rect 303 -956 307 -949
rect 303 -968 307 -961
rect 226 -990 230 -976
rect 242 -990 246 -976
rect 280 -990 284 -976
rect 300 -990 304 -976
rect 226 -994 311 -990
rect 373 -999 378 -945
rect 568 -948 576 -946
rect 516 -952 576 -948
rect 522 -964 526 -952
rect 550 -964 554 -952
rect 568 -954 576 -952
rect 498 -983 523 -979
rect 410 -990 475 -986
rect 540 -984 544 -970
rect 558 -984 562 -970
rect 482 -990 505 -986
rect 512 -990 533 -986
rect 540 -988 551 -984
rect 558 -988 573 -984
rect 410 -991 415 -990
rect 540 -994 544 -988
rect 531 -998 544 -994
rect 218 -1004 310 -1000
rect 218 -1008 230 -1004
rect 226 -1017 230 -1008
rect 242 -1017 246 -1004
rect 280 -1017 284 -1004
rect 300 -1017 304 -1004
rect 373 -1005 423 -999
rect 431 -1005 482 -999
rect 531 -1002 535 -998
rect 558 -1002 562 -988
rect 522 -1013 526 -1006
rect 540 -1013 544 -1006
rect 586 -1005 592 -942
rect 707 -940 718 -938
rect 775 -940 779 -933
rect 906 -936 993 -932
rect 1080 -933 1086 -931
rect 1105 -933 1109 -914
rect 1132 -924 1136 -914
rect 906 -940 918 -936
rect 707 -944 794 -940
rect 914 -951 918 -940
rect 933 -951 937 -936
rect 953 -951 957 -936
rect 975 -951 979 -936
rect 1080 -937 1098 -933
rect 1105 -937 1124 -933
rect 1080 -945 1091 -941
rect 1080 -948 1087 -945
rect 1105 -956 1109 -937
rect 1132 -956 1136 -929
rect 1163 -933 1167 -914
rect 1326 -925 1330 -916
rect 1338 -925 1342 -822
rect 1360 -822 1364 -815
rect 1374 -822 1394 -818
rect 1364 -835 1366 -831
rect 1364 -836 1369 -835
rect 1198 -929 1279 -925
rect 1310 -928 1342 -925
rect 1348 -926 1352 -916
rect 1374 -926 1378 -822
rect 1398 -822 1402 -815
rect 1386 -834 1390 -831
rect 1413 -834 1509 -829
rect 1381 -835 1390 -834
rect 1386 -836 1390 -835
rect 1416 -838 1420 -834
rect 1503 -862 1509 -834
rect 1503 -866 1528 -862
rect 1510 -870 1514 -866
rect 1398 -885 1406 -883
rect 1398 -886 1417 -885
rect 1402 -889 1417 -886
rect 1424 -886 1428 -878
rect 1518 -886 1522 -878
rect 1402 -901 1406 -889
rect 1424 -890 1511 -886
rect 1518 -890 1531 -886
rect 1424 -892 1428 -890
rect 1310 -931 1314 -928
rect 1348 -931 1378 -926
rect 1154 -937 1167 -933
rect 1163 -956 1167 -937
rect 1174 -940 1178 -933
rect 1174 -952 1178 -945
rect 859 -965 866 -962
rect 923 -965 927 -957
rect 943 -965 947 -957
rect 983 -965 987 -957
rect 859 -969 915 -965
rect 923 -969 976 -965
rect 983 -969 1004 -965
rect 706 -976 785 -972
rect 853 -976 925 -972
rect 706 -980 718 -976
rect 714 -991 718 -980
rect 733 -991 737 -976
rect 767 -991 771 -976
rect 817 -979 824 -976
rect 817 -983 935 -979
rect 835 -990 945 -986
rect 835 -991 841 -990
rect 953 -994 957 -969
rect 983 -994 987 -969
rect 999 -970 1004 -969
rect 1097 -970 1101 -960
rect 1089 -974 1101 -970
rect 1113 -974 1117 -960
rect 1151 -974 1155 -960
rect 1171 -974 1175 -960
rect 1089 -978 1182 -974
rect 1318 -983 1322 -951
rect 1348 -934 1352 -931
rect 1364 -976 1368 -974
rect 1518 -893 1522 -890
rect 1510 -901 1514 -897
rect 1503 -905 1528 -901
rect 1416 -921 1420 -912
rect 1503 -921 1507 -905
rect 1410 -925 1507 -921
rect 1386 -947 1390 -941
rect 1410 -947 1413 -925
rect 1386 -951 1413 -947
rect 1386 -976 1390 -951
rect 1364 -980 1390 -976
rect 1364 -983 1368 -980
rect 1318 -987 1368 -983
rect 723 -1005 727 -997
rect 743 -1005 747 -997
rect 775 -1005 779 -997
rect 1097 -993 1312 -989
rect 914 -1005 918 -998
rect 975 -1005 979 -998
rect 989 -1005 997 -1002
rect 550 -1013 554 -1006
rect 586 -1009 715 -1005
rect 723 -1009 768 -1005
rect 775 -1009 805 -1005
rect 907 -1009 997 -1005
rect 1097 -1006 1101 -993
rect 1113 -1006 1117 -993
rect 1151 -1006 1155 -993
rect 1171 -1006 1175 -993
rect 570 -1013 576 -1010
rect 515 -1017 576 -1013
rect 620 -1016 725 -1012
rect 620 -1019 626 -1016
rect 475 -1022 482 -1020
rect 620 -1022 625 -1019
rect 53 -1042 141 -1039
rect 234 -1042 238 -1023
rect 261 -1033 265 -1023
rect 53 -1046 227 -1042
rect 234 -1046 253 -1042
rect -17 -1232 -13 -1220
rect 5 -1221 39 -1217
rect 47 -1054 220 -1049
rect 5 -1223 9 -1221
rect -109 -1262 -105 -1259
rect -71 -1262 -41 -1257
rect -235 -1307 -231 -1282
rect -257 -1311 -231 -1307
rect -257 -1314 -253 -1311
rect -303 -1318 -253 -1314
rect -101 -1314 -97 -1282
rect -71 -1265 -67 -1262
rect -55 -1307 -51 -1305
rect -3 -1252 1 -1243
rect -9 -1256 7 -1252
rect -33 -1278 -29 -1272
rect -9 -1278 -6 -1256
rect -33 -1282 -6 -1278
rect -33 -1307 -29 -1282
rect -55 -1311 -29 -1307
rect -55 -1314 -51 -1311
rect -101 -1318 -51 -1314
rect -299 -1330 -219 -1326
rect -307 -1337 -303 -1333
rect -299 -1337 -295 -1330
rect -283 -1337 -265 -1333
rect -308 -1350 -307 -1344
rect -311 -1351 -307 -1350
rect -295 -1440 -291 -1431
rect -283 -1440 -279 -1337
rect -261 -1337 -257 -1330
rect -247 -1337 -227 -1333
rect -257 -1350 -255 -1346
rect -257 -1351 -252 -1350
rect -311 -1443 -279 -1440
rect -273 -1441 -269 -1431
rect -247 -1441 -243 -1337
rect -223 -1337 -219 -1330
rect -94 -1328 -14 -1324
rect -102 -1335 -98 -1331
rect -94 -1335 -90 -1328
rect -78 -1335 -60 -1331
rect -235 -1349 -231 -1346
rect -208 -1349 -187 -1344
rect -103 -1348 -102 -1342
rect -106 -1349 -102 -1348
rect -240 -1350 -231 -1349
rect -235 -1351 -231 -1350
rect -205 -1353 -201 -1349
rect -223 -1400 -215 -1398
rect -223 -1401 -204 -1400
rect -219 -1404 -204 -1401
rect -197 -1401 -193 -1393
rect -219 -1416 -215 -1404
rect -197 -1405 -176 -1401
rect -197 -1407 -193 -1405
rect -311 -1446 -307 -1443
rect -273 -1446 -243 -1441
rect -303 -1498 -299 -1466
rect -273 -1449 -269 -1446
rect -257 -1491 -253 -1489
rect -205 -1436 -201 -1427
rect -211 -1440 -187 -1436
rect -90 -1438 -86 -1429
rect -78 -1438 -74 -1335
rect -56 -1335 -52 -1328
rect -42 -1335 -22 -1331
rect -52 -1348 -50 -1344
rect -52 -1349 -47 -1348
rect -235 -1462 -231 -1456
rect -211 -1462 -208 -1440
rect -235 -1466 -208 -1462
rect -106 -1441 -74 -1438
rect -68 -1439 -64 -1429
rect -42 -1439 -38 -1335
rect -18 -1335 -14 -1328
rect -30 -1347 -26 -1344
rect -3 -1347 18 -1342
rect -35 -1348 -26 -1347
rect -30 -1349 -26 -1348
rect 0 -1351 4 -1347
rect -18 -1398 -10 -1396
rect -18 -1399 1 -1398
rect -14 -1402 1 -1399
rect 8 -1399 12 -1391
rect 47 -1399 58 -1054
rect 78 -1057 85 -1054
rect 234 -1065 238 -1046
rect 261 -1065 265 -1038
rect 292 -1042 296 -1023
rect 475 -1027 625 -1022
rect 632 -1023 735 -1019
rect 632 -1025 639 -1023
rect 743 -1026 747 -1009
rect 775 -1026 779 -1009
rect 800 -1010 805 -1009
rect 1320 -1004 1400 -1000
rect 1287 -1011 1316 -1007
rect 327 -1038 406 -1033
rect 521 -1035 601 -1031
rect 283 -1046 296 -1042
rect 292 -1065 296 -1046
rect 303 -1049 307 -1042
rect 303 -1061 307 -1054
rect 527 -1050 531 -1035
rect 546 -1050 550 -1035
rect 580 -1050 584 -1035
rect 593 -1039 601 -1035
rect 619 -1041 625 -1027
rect 714 -1035 718 -1030
rect 707 -1037 718 -1035
rect 767 -1037 771 -1030
rect 1020 -1031 1028 -1027
rect 1105 -1031 1109 -1012
rect 1132 -1022 1136 -1012
rect 906 -1037 985 -1033
rect 1020 -1035 1098 -1031
rect 1105 -1035 1124 -1031
rect 707 -1041 786 -1037
rect 906 -1041 918 -1037
rect 536 -1064 540 -1056
rect 556 -1064 560 -1056
rect 588 -1064 592 -1056
rect 914 -1052 918 -1041
rect 933 -1052 937 -1037
rect 967 -1052 971 -1037
rect 1081 -1043 1091 -1039
rect 1105 -1054 1109 -1035
rect 1132 -1054 1136 -1027
rect 1163 -1031 1167 -1012
rect 1198 -1027 1281 -1023
rect 1154 -1035 1167 -1031
rect 1163 -1054 1167 -1035
rect 1174 -1038 1178 -1031
rect 1174 -1050 1178 -1043
rect 498 -1068 528 -1064
rect 536 -1068 581 -1064
rect 588 -1068 610 -1064
rect 705 -1067 774 -1063
rect 923 -1066 927 -1058
rect 943 -1066 947 -1058
rect 975 -1066 979 -1058
rect 226 -1079 230 -1069
rect 227 -1083 230 -1079
rect 242 -1083 246 -1069
rect 280 -1083 284 -1069
rect 300 -1083 304 -1069
rect 486 -1071 492 -1069
rect 486 -1075 538 -1071
rect 475 -1078 482 -1076
rect 475 -1082 548 -1078
rect 475 -1083 482 -1082
rect 227 -1087 311 -1083
rect 556 -1085 560 -1068
rect 588 -1085 592 -1068
rect 705 -1071 717 -1067
rect 713 -1082 717 -1071
rect 732 -1082 736 -1067
rect 756 -1082 760 -1067
rect 812 -1070 915 -1066
rect 923 -1070 968 -1066
rect 975 -1070 999 -1066
rect 1097 -1068 1101 -1058
rect 817 -1077 925 -1073
rect 817 -1079 824 -1077
rect 835 -1084 935 -1080
rect 835 -1085 841 -1084
rect 943 -1087 947 -1070
rect 975 -1087 979 -1070
rect 993 -1072 999 -1070
rect 1089 -1072 1101 -1068
rect 1113 -1072 1117 -1058
rect 1151 -1072 1155 -1058
rect 1171 -1072 1175 -1058
rect 1089 -1076 1182 -1072
rect 1213 -1081 1220 -1079
rect 1213 -1085 1226 -1081
rect 273 -1096 415 -1091
rect 527 -1096 531 -1089
rect 580 -1096 584 -1089
rect 594 -1096 600 -1093
rect 722 -1096 726 -1088
rect 764 -1096 768 -1088
rect 520 -1100 600 -1096
rect 649 -1100 714 -1096
rect 722 -1100 757 -1096
rect 764 -1100 778 -1096
rect 914 -1098 918 -1091
rect 967 -1098 971 -1091
rect 1091 -1093 1181 -1089
rect 980 -1098 988 -1095
rect 1091 -1098 1101 -1093
rect 227 -1106 297 -1102
rect 227 -1111 240 -1106
rect 236 -1121 240 -1111
rect 255 -1121 259 -1106
rect 279 -1121 283 -1106
rect 632 -1109 724 -1105
rect 732 -1114 736 -1100
rect 764 -1114 768 -1100
rect 907 -1102 988 -1098
rect 1097 -1106 1101 -1098
rect 1113 -1106 1117 -1093
rect 1151 -1106 1155 -1093
rect 1171 -1106 1175 -1093
rect 521 -1121 592 -1117
rect 245 -1135 249 -1127
rect 287 -1135 291 -1127
rect 225 -1139 237 -1135
rect 245 -1139 280 -1135
rect 287 -1139 354 -1135
rect 225 -1140 230 -1139
rect 225 -1148 247 -1144
rect 225 -1151 232 -1148
rect 255 -1153 259 -1139
rect 287 -1153 291 -1139
rect 349 -1142 354 -1139
rect 527 -1136 531 -1121
rect 546 -1136 550 -1121
rect 570 -1136 574 -1121
rect 584 -1125 592 -1121
rect 713 -1123 717 -1118
rect 706 -1125 717 -1123
rect 756 -1125 760 -1118
rect 904 -1124 973 -1120
rect 706 -1129 773 -1125
rect 904 -1128 916 -1124
rect 475 -1150 482 -1148
rect 536 -1150 540 -1142
rect 578 -1150 582 -1142
rect 912 -1139 916 -1128
rect 931 -1139 935 -1124
rect 955 -1139 959 -1124
rect 1105 -1131 1109 -1112
rect 1132 -1122 1136 -1112
rect 1040 -1135 1098 -1131
rect 1105 -1135 1124 -1131
rect 1028 -1143 1091 -1139
rect 703 -1149 782 -1145
rect 475 -1155 528 -1150
rect 536 -1154 571 -1150
rect 578 -1154 610 -1150
rect 703 -1153 715 -1149
rect 236 -1160 240 -1157
rect 229 -1164 240 -1160
rect 279 -1164 283 -1157
rect 464 -1159 471 -1156
rect 464 -1163 538 -1159
rect 229 -1168 298 -1164
rect 546 -1168 550 -1154
rect 578 -1168 582 -1154
rect 711 -1161 715 -1153
rect 759 -1161 763 -1149
rect 921 -1153 925 -1145
rect 963 -1153 967 -1145
rect 797 -1157 913 -1153
rect 921 -1157 956 -1153
rect 963 -1157 993 -1153
rect 1105 -1154 1109 -1135
rect 1132 -1154 1136 -1127
rect 1163 -1131 1167 -1112
rect 1287 -1123 1293 -1011
rect 1320 -1011 1324 -1004
rect 1336 -1011 1354 -1007
rect 1311 -1024 1312 -1018
rect 1308 -1025 1312 -1024
rect 1324 -1114 1328 -1105
rect 1336 -1114 1340 -1011
rect 1358 -1011 1362 -1004
rect 1372 -1011 1392 -1007
rect 1362 -1024 1364 -1020
rect 1362 -1025 1367 -1024
rect 1198 -1127 1293 -1123
rect 1308 -1117 1340 -1114
rect 1346 -1115 1350 -1105
rect 1372 -1115 1376 -1011
rect 1396 -1011 1400 -1004
rect 1384 -1023 1388 -1020
rect 1411 -1023 1507 -1018
rect 1379 -1024 1388 -1023
rect 1384 -1025 1388 -1024
rect 1414 -1027 1418 -1023
rect 1502 -1051 1507 -1023
rect 1502 -1055 1527 -1051
rect 1509 -1059 1513 -1055
rect 1396 -1074 1404 -1072
rect 1396 -1075 1415 -1074
rect 1400 -1078 1415 -1075
rect 1422 -1075 1426 -1067
rect 1517 -1075 1521 -1067
rect 1400 -1090 1404 -1078
rect 1422 -1079 1510 -1075
rect 1517 -1079 1530 -1075
rect 1422 -1081 1426 -1079
rect 1308 -1120 1312 -1117
rect 1346 -1120 1376 -1115
rect 1154 -1135 1167 -1131
rect 1163 -1154 1167 -1135
rect 1174 -1138 1178 -1131
rect 1174 -1150 1178 -1143
rect 226 -1181 296 -1177
rect 527 -1179 531 -1172
rect 570 -1179 574 -1172
rect 691 -1176 696 -1175
rect 585 -1179 591 -1176
rect 226 -1186 239 -1181
rect 235 -1196 239 -1186
rect 254 -1196 258 -1181
rect 278 -1196 282 -1181
rect 520 -1183 591 -1179
rect 691 -1180 712 -1176
rect 749 -1181 753 -1167
rect 767 -1181 771 -1167
rect 682 -1183 687 -1182
rect 682 -1187 722 -1183
rect 749 -1185 760 -1181
rect 767 -1185 791 -1181
rect 669 -1190 675 -1188
rect 669 -1194 732 -1190
rect 584 -1199 592 -1197
rect 224 -1210 229 -1209
rect 244 -1210 248 -1202
rect 286 -1210 290 -1202
rect 520 -1203 592 -1199
rect 224 -1214 236 -1210
rect 244 -1214 279 -1210
rect 286 -1214 372 -1210
rect 224 -1223 246 -1219
rect 224 -1226 231 -1223
rect 254 -1228 258 -1214
rect 286 -1228 290 -1214
rect 367 -1215 372 -1214
rect 526 -1215 530 -1203
rect 564 -1215 568 -1203
rect 584 -1205 592 -1203
rect 624 -1201 741 -1197
rect 512 -1230 518 -1228
rect 235 -1235 239 -1232
rect 228 -1239 239 -1235
rect 278 -1239 282 -1232
rect 512 -1234 527 -1230
rect 554 -1235 558 -1221
rect 572 -1235 576 -1221
rect 607 -1235 613 -1234
rect 228 -1243 297 -1239
rect 502 -1241 537 -1237
rect 554 -1239 565 -1235
rect 572 -1239 613 -1235
rect 411 -1245 547 -1244
rect 411 -1248 502 -1245
rect 226 -1256 296 -1252
rect 226 -1261 239 -1256
rect 235 -1271 239 -1261
rect 254 -1271 258 -1256
rect 278 -1271 282 -1256
rect 224 -1285 229 -1284
rect 244 -1285 248 -1277
rect 286 -1285 290 -1277
rect 411 -1281 417 -1248
rect 508 -1248 547 -1245
rect 554 -1252 558 -1239
rect 535 -1256 558 -1252
rect 535 -1260 539 -1256
rect 554 -1260 558 -1256
rect 572 -1260 576 -1239
rect 526 -1270 530 -1264
rect 519 -1271 530 -1270
rect 544 -1271 548 -1264
rect 564 -1271 568 -1264
rect 582 -1271 588 -1268
rect 519 -1275 588 -1271
rect 519 -1277 526 -1275
rect 337 -1285 417 -1281
rect 224 -1289 236 -1285
rect 244 -1289 279 -1285
rect 286 -1289 343 -1285
rect 624 -1288 629 -1201
rect 749 -1205 753 -1185
rect 720 -1209 753 -1205
rect 720 -1213 724 -1209
rect 739 -1213 743 -1209
rect 767 -1213 771 -1185
rect 784 -1186 791 -1185
rect 711 -1222 715 -1217
rect 704 -1224 715 -1222
rect 729 -1224 733 -1217
rect 749 -1224 753 -1217
rect 759 -1224 763 -1217
rect 704 -1228 782 -1224
rect 797 -1288 803 -1157
rect 835 -1166 923 -1162
rect 835 -1167 841 -1166
rect 931 -1171 935 -1157
rect 963 -1171 967 -1157
rect 987 -1159 993 -1157
rect 1097 -1168 1101 -1158
rect 1089 -1172 1101 -1168
rect 1113 -1172 1117 -1158
rect 1151 -1172 1155 -1158
rect 1171 -1172 1175 -1158
rect 1316 -1172 1320 -1140
rect 1346 -1123 1350 -1120
rect 1362 -1165 1366 -1163
rect 1517 -1082 1521 -1079
rect 1509 -1090 1513 -1086
rect 1502 -1094 1527 -1090
rect 1414 -1110 1418 -1101
rect 1502 -1110 1507 -1094
rect 1408 -1114 1507 -1110
rect 1384 -1136 1388 -1130
rect 1408 -1136 1411 -1114
rect 1384 -1140 1411 -1136
rect 1384 -1165 1388 -1140
rect 1362 -1169 1388 -1165
rect 1362 -1172 1366 -1169
rect 912 -1182 916 -1175
rect 955 -1182 959 -1175
rect 1089 -1176 1182 -1172
rect 1316 -1176 1366 -1172
rect 967 -1182 974 -1180
rect 905 -1186 974 -1182
rect 1086 -1191 1181 -1187
rect 1086 -1194 1102 -1191
rect 1086 -1196 1101 -1194
rect 1097 -1204 1101 -1196
rect 1113 -1204 1117 -1191
rect 1151 -1204 1155 -1191
rect 1171 -1204 1175 -1191
rect 1321 -1193 1401 -1189
rect 1266 -1197 1317 -1193
rect 903 -1218 991 -1214
rect 903 -1222 915 -1218
rect 911 -1230 915 -1222
rect 968 -1230 972 -1218
rect 1105 -1229 1109 -1210
rect 1132 -1220 1136 -1210
rect 1061 -1233 1098 -1229
rect 1105 -1233 1124 -1229
rect 1061 -1235 1067 -1233
rect 896 -1249 912 -1245
rect 959 -1250 963 -1236
rect 976 -1250 980 -1236
rect 1077 -1237 1083 -1236
rect 1077 -1241 1091 -1237
rect 885 -1256 922 -1252
rect 959 -1254 969 -1250
rect 976 -1254 1001 -1250
rect 1105 -1252 1109 -1233
rect 1132 -1252 1136 -1225
rect 1163 -1229 1167 -1210
rect 1266 -1221 1271 -1197
rect 1313 -1200 1317 -1197
rect 1321 -1200 1325 -1193
rect 1337 -1200 1355 -1196
rect 1312 -1213 1313 -1207
rect 1198 -1225 1271 -1221
rect 1309 -1214 1313 -1213
rect 1154 -1233 1167 -1229
rect 1163 -1252 1167 -1233
rect 1174 -1236 1178 -1229
rect 1174 -1248 1178 -1241
rect 875 -1263 932 -1259
rect 865 -1270 941 -1266
rect 224 -1298 246 -1294
rect 224 -1301 231 -1298
rect 254 -1303 258 -1289
rect 286 -1303 290 -1289
rect 367 -1294 803 -1288
rect 859 -1277 951 -1273
rect 235 -1310 239 -1307
rect 228 -1314 239 -1310
rect 278 -1314 282 -1307
rect 358 -1310 824 -1303
rect 228 -1318 297 -1314
rect 337 -1325 841 -1319
rect 226 -1331 296 -1327
rect 226 -1336 239 -1331
rect 235 -1346 239 -1336
rect 254 -1346 258 -1331
rect 278 -1346 282 -1331
rect 859 -1333 866 -1277
rect 959 -1281 963 -1254
rect 920 -1285 963 -1281
rect 920 -1289 924 -1285
rect 939 -1289 943 -1285
rect 959 -1289 963 -1285
rect 976 -1289 980 -1254
rect 1097 -1266 1101 -1256
rect 1089 -1270 1101 -1266
rect 1113 -1270 1117 -1256
rect 1151 -1270 1155 -1256
rect 1171 -1270 1175 -1256
rect 1089 -1274 1182 -1270
rect 911 -1299 915 -1293
rect 904 -1300 915 -1299
rect 929 -1300 933 -1293
rect 949 -1300 953 -1293
rect 968 -1300 972 -1293
rect 984 -1300 991 -1298
rect 904 -1301 991 -1300
rect 1097 -1301 1101 -1274
rect 904 -1304 1101 -1301
rect 1325 -1303 1329 -1294
rect 1337 -1303 1341 -1200
rect 1359 -1200 1363 -1193
rect 1373 -1200 1393 -1196
rect 1363 -1213 1365 -1209
rect 1363 -1214 1368 -1213
rect 904 -1305 911 -1304
rect 1309 -1306 1341 -1303
rect 1347 -1304 1351 -1294
rect 1373 -1304 1377 -1200
rect 1397 -1200 1401 -1193
rect 1385 -1212 1389 -1209
rect 1412 -1212 1507 -1207
rect 1380 -1213 1389 -1212
rect 1385 -1214 1389 -1213
rect 1415 -1216 1419 -1212
rect 1499 -1213 1507 -1212
rect 1500 -1240 1507 -1213
rect 1500 -1244 1525 -1240
rect 1507 -1248 1511 -1244
rect 1397 -1263 1405 -1261
rect 1397 -1264 1416 -1263
rect 1401 -1267 1416 -1264
rect 1423 -1264 1427 -1256
rect 1515 -1264 1519 -1256
rect 1401 -1279 1405 -1267
rect 1423 -1268 1508 -1264
rect 1515 -1268 1528 -1264
rect 1423 -1270 1427 -1268
rect 1309 -1309 1313 -1306
rect 1347 -1309 1377 -1304
rect 926 -1311 936 -1310
rect 926 -1317 1083 -1311
rect 926 -1318 936 -1317
rect 349 -1339 866 -1333
rect 224 -1360 229 -1359
rect 244 -1360 248 -1352
rect 286 -1360 290 -1352
rect 386 -1360 391 -1359
rect 224 -1364 236 -1360
rect 244 -1364 279 -1360
rect 286 -1364 391 -1360
rect 224 -1373 246 -1369
rect 224 -1376 231 -1373
rect 254 -1378 258 -1364
rect 286 -1378 290 -1364
rect 235 -1385 239 -1382
rect 228 -1389 239 -1385
rect 278 -1389 282 -1382
rect 228 -1393 297 -1389
rect -14 -1414 -10 -1402
rect 8 -1403 58 -1399
rect 8 -1405 12 -1403
rect -106 -1444 -102 -1441
rect -68 -1444 -38 -1439
rect -235 -1491 -231 -1466
rect -257 -1495 -231 -1491
rect -257 -1498 -253 -1495
rect -303 -1502 -253 -1498
rect -98 -1496 -94 -1464
rect -68 -1447 -64 -1444
rect -52 -1489 -48 -1487
rect 607 -1408 613 -1360
rect 659 -1387 665 -1362
rect 785 -1375 792 -1355
rect 785 -1383 793 -1375
rect 996 -1377 1001 -1345
rect 1046 -1351 1062 -1334
rect 659 -1388 1013 -1387
rect 659 -1394 1014 -1388
rect 1050 -1408 1059 -1351
rect 1317 -1361 1321 -1329
rect 1347 -1312 1351 -1309
rect 1363 -1354 1367 -1352
rect 1515 -1271 1519 -1268
rect 1507 -1279 1511 -1275
rect 1500 -1283 1525 -1279
rect 1415 -1299 1419 -1290
rect 1500 -1299 1503 -1283
rect 1409 -1303 1503 -1299
rect 1385 -1325 1389 -1319
rect 1409 -1325 1412 -1303
rect 1385 -1329 1412 -1325
rect 1385 -1354 1389 -1329
rect 1363 -1358 1389 -1354
rect 1363 -1361 1367 -1358
rect 1317 -1365 1367 -1361
rect 1322 -1381 1402 -1377
rect 1314 -1388 1318 -1384
rect 1322 -1388 1326 -1381
rect 1338 -1388 1356 -1384
rect 1313 -1401 1314 -1395
rect 607 -1415 1059 -1408
rect 1310 -1402 1314 -1401
rect 0 -1434 4 -1425
rect -6 -1438 18 -1434
rect -30 -1460 -26 -1454
rect -6 -1460 -3 -1438
rect -30 -1464 -3 -1460
rect -30 -1489 -26 -1464
rect -52 -1493 -26 -1489
rect 1326 -1491 1330 -1482
rect 1338 -1491 1342 -1388
rect 1360 -1388 1364 -1381
rect 1374 -1388 1394 -1384
rect 1364 -1401 1366 -1397
rect 1364 -1402 1369 -1401
rect -52 -1496 -48 -1493
rect -98 -1500 -48 -1496
rect 1310 -1494 1342 -1491
rect 1348 -1492 1352 -1482
rect 1374 -1492 1378 -1388
rect 1398 -1388 1402 -1381
rect 1386 -1400 1390 -1397
rect 1413 -1400 1510 -1395
rect 1381 -1401 1390 -1400
rect 1386 -1402 1390 -1401
rect 1416 -1404 1420 -1400
rect 1503 -1428 1510 -1400
rect 1503 -1432 1528 -1428
rect 1510 -1436 1514 -1432
rect 1398 -1451 1406 -1449
rect 1398 -1452 1417 -1451
rect 1402 -1455 1417 -1452
rect 1424 -1452 1428 -1444
rect 1518 -1452 1522 -1444
rect 1402 -1467 1406 -1455
rect 1424 -1456 1511 -1452
rect 1518 -1456 1531 -1452
rect 1424 -1458 1428 -1456
rect 1310 -1497 1314 -1494
rect 1348 -1497 1378 -1492
rect 1318 -1549 1322 -1517
rect 1348 -1500 1352 -1497
rect 1364 -1542 1368 -1540
rect 1518 -1459 1522 -1456
rect 1510 -1467 1514 -1463
rect 1503 -1471 1528 -1467
rect 1416 -1487 1420 -1478
rect 1503 -1487 1507 -1471
rect 1410 -1491 1507 -1487
rect 1386 -1513 1390 -1507
rect 1410 -1513 1413 -1491
rect 1386 -1517 1413 -1513
rect 1386 -1542 1390 -1517
rect 1364 -1546 1390 -1542
rect 1364 -1549 1368 -1546
rect 1318 -1553 1368 -1549
<< m2contact >>
rect 1305 -645 1310 -639
rect -311 -781 -306 -775
rect -253 -781 -248 -776
rect 261 -761 266 -756
rect -238 -780 -233 -774
rect -212 -780 -206 -774
rect 220 -777 225 -772
rect -116 -801 -111 -795
rect -58 -801 -53 -796
rect -43 -800 -38 -794
rect -17 -800 -11 -794
rect 322 -761 327 -756
rect 302 -777 307 -772
rect -313 -972 -308 -966
rect -255 -972 -250 -967
rect 261 -853 266 -848
rect 220 -869 225 -864
rect -240 -971 -235 -965
rect -214 -971 -208 -965
rect -115 -984 -110 -978
rect -57 -984 -52 -979
rect -42 -983 -37 -977
rect -16 -983 -10 -977
rect 322 -853 327 -848
rect 1363 -645 1368 -640
rect 1378 -644 1383 -638
rect 1404 -644 1410 -638
rect 302 -869 307 -864
rect 1308 -835 1313 -829
rect 475 -882 482 -877
rect 848 -877 853 -872
rect 636 -904 642 -899
rect 261 -945 266 -940
rect 220 -961 225 -956
rect -313 -1166 -308 -1160
rect -255 -1166 -250 -1161
rect -240 -1165 -235 -1159
rect -214 -1165 -208 -1159
rect -111 -1166 -106 -1160
rect -53 -1166 -48 -1161
rect -38 -1165 -33 -1159
rect -12 -1165 -6 -1159
rect 322 -945 327 -940
rect 302 -961 307 -956
rect 475 -990 482 -983
rect 573 -988 579 -982
rect 423 -1005 431 -999
rect 1132 -929 1137 -924
rect 1091 -945 1096 -940
rect 1193 -929 1198 -924
rect 1366 -835 1371 -830
rect 1381 -834 1386 -828
rect 1407 -834 1413 -828
rect 1173 -945 1178 -940
rect 848 -976 853 -971
rect 261 -1038 266 -1033
rect 220 -1054 225 -1049
rect -313 -1350 -308 -1344
rect -255 -1350 -250 -1345
rect -240 -1349 -235 -1343
rect -214 -1349 -208 -1343
rect -108 -1348 -103 -1342
rect -50 -1348 -45 -1343
rect -35 -1347 -30 -1341
rect -9 -1347 -3 -1341
rect 322 -1038 327 -1033
rect 302 -1054 307 -1049
rect 1132 -1027 1137 -1022
rect 619 -1049 625 -1041
rect 1091 -1043 1096 -1038
rect 1193 -1027 1198 -1022
rect 1173 -1043 1178 -1038
rect 807 -1071 812 -1066
rect 643 -1101 649 -1096
rect 1032 -1135 1040 -1130
rect 1132 -1127 1137 -1122
rect 1091 -1143 1096 -1138
rect 1193 -1127 1198 -1122
rect 1306 -1024 1311 -1018
rect 1364 -1024 1369 -1019
rect 1379 -1023 1384 -1017
rect 1405 -1023 1411 -1017
rect 1173 -1143 1178 -1138
rect 502 -1251 508 -1245
rect 643 -1283 649 -1276
rect 1132 -1225 1137 -1220
rect 1091 -1241 1096 -1236
rect 1193 -1225 1198 -1220
rect 1307 -1213 1312 -1207
rect 1173 -1241 1178 -1236
rect 1365 -1213 1370 -1208
rect 1380 -1212 1385 -1206
rect 1406 -1212 1412 -1206
rect 1308 -1401 1313 -1395
rect 1366 -1401 1371 -1396
rect 1381 -1400 1386 -1394
rect 1407 -1400 1413 -1394
<< metal2 >>
rect 1310 -640 1378 -639
rect 1310 -643 1363 -640
rect 1368 -643 1378 -640
rect 1383 -643 1404 -639
rect 266 -761 322 -757
rect -306 -776 -238 -775
rect -306 -779 -253 -776
rect -248 -779 -238 -776
rect -233 -779 -212 -775
rect 225 -777 302 -772
rect -111 -796 -43 -795
rect -111 -799 -58 -796
rect -53 -799 -43 -796
rect -38 -799 -17 -795
rect 475 -803 895 -796
rect 266 -853 322 -849
rect -184 -861 31 -855
rect -308 -967 -240 -966
rect -308 -970 -255 -967
rect -250 -970 -240 -967
rect -235 -970 -214 -966
rect -184 -1028 -176 -861
rect 225 -869 302 -864
rect 475 -877 482 -803
rect 266 -945 322 -941
rect -172 -953 60 -945
rect -172 -954 52 -953
rect -172 -1047 -160 -954
rect 225 -961 302 -956
rect -110 -979 -42 -978
rect -110 -982 -57 -979
rect -52 -982 -42 -979
rect -37 -982 -16 -978
rect 475 -983 482 -882
rect 636 -899 642 -803
rect 889 -855 895 -803
rect 1313 -830 1381 -829
rect 1313 -833 1366 -830
rect 1371 -833 1381 -830
rect 1386 -833 1407 -829
rect 848 -971 853 -877
rect 1137 -929 1193 -925
rect 1096 -945 1173 -940
rect 579 -988 662 -982
rect 266 -1038 322 -1034
rect -184 -1058 -160 -1047
rect -308 -1161 -240 -1160
rect -308 -1164 -255 -1161
rect -250 -1164 -240 -1161
rect -235 -1164 -214 -1160
rect -184 -1221 -177 -1058
rect -106 -1161 -38 -1160
rect -106 -1164 -53 -1161
rect -48 -1164 -38 -1161
rect -33 -1164 -12 -1160
rect -308 -1345 -240 -1344
rect -308 -1348 -255 -1345
rect -250 -1348 -240 -1345
rect -235 -1348 -214 -1344
rect -103 -1343 -35 -1342
rect -103 -1346 -50 -1343
rect -45 -1346 -35 -1343
rect -30 -1346 -9 -1342
rect 53 -1398 70 -1039
rect 225 -1054 302 -1049
rect -183 -1409 70 -1398
rect 423 -1397 431 -1005
rect 848 -1044 853 -976
rect 1137 -1027 1193 -1023
rect 1311 -1019 1379 -1018
rect 1311 -1022 1364 -1019
rect 1369 -1022 1379 -1019
rect 1384 -1022 1405 -1018
rect 1096 -1043 1173 -1038
rect 625 -1049 853 -1044
rect 502 -1278 508 -1251
rect 643 -1276 649 -1101
rect 502 -1283 643 -1278
rect 807 -1278 812 -1071
rect 1137 -1127 1193 -1123
rect 649 -1283 812 -1278
rect 1032 -1397 1040 -1135
rect 1096 -1143 1173 -1138
rect 1312 -1208 1380 -1207
rect 1312 -1211 1365 -1208
rect 1370 -1211 1380 -1208
rect 1385 -1211 1406 -1207
rect 1137 -1225 1193 -1221
rect 1096 -1241 1173 -1236
rect 423 -1405 1040 -1397
rect 1313 -1396 1381 -1395
rect 1313 -1399 1366 -1396
rect 1371 -1399 1381 -1396
rect 1386 -1399 1407 -1395
rect 53 -1410 70 -1409
<< m3contact >>
rect 337 -761 343 -756
rect 112 -779 119 -772
rect 358 -853 364 -848
rect 101 -871 108 -864
rect 619 -828 627 -821
rect 386 -884 391 -879
rect 464 -885 471 -879
rect 400 -893 405 -888
rect 464 -942 471 -935
rect 89 -963 96 -956
rect 594 -888 603 -879
rect 486 -893 492 -888
rect 1011 -864 1016 -859
rect 817 -886 824 -880
rect 835 -893 841 -888
rect 620 -910 626 -903
rect 801 -905 806 -900
rect 620 -920 626 -914
rect 632 -926 639 -921
rect 859 -969 866 -962
rect 999 -970 1004 -965
rect 498 -981 505 -975
rect 410 -991 415 -986
rect 498 -994 505 -987
rect 817 -983 824 -976
rect 835 -991 841 -986
rect 475 -1005 482 -999
rect 400 -1038 405 -1033
rect 78 -1057 85 -1049
rect 273 -1096 278 -1091
rect 410 -1096 415 -1091
rect 349 -1142 354 -1135
rect 225 -1151 232 -1144
rect 367 -1215 372 -1210
rect 224 -1226 231 -1219
rect 367 -1294 372 -1288
rect 224 -1301 231 -1294
rect 358 -1310 363 -1303
rect 337 -1325 343 -1319
rect 349 -1339 354 -1333
rect 386 -1364 391 -1359
rect 224 -1376 231 -1369
rect 800 -1010 805 -1005
rect 620 -1019 626 -1012
rect 475 -1027 482 -1020
rect 632 -1025 639 -1019
rect 498 -1068 505 -1062
rect 486 -1075 492 -1069
rect 604 -1070 610 -1064
rect 475 -1083 482 -1076
rect 632 -1111 639 -1105
rect 475 -1155 482 -1148
rect 604 -1156 610 -1150
rect 464 -1163 471 -1156
rect 512 -1234 518 -1228
rect 502 -1241 508 -1235
rect 691 -1180 696 -1175
rect 682 -1187 687 -1182
rect 669 -1194 675 -1188
rect 993 -1072 999 -1066
rect 817 -1079 824 -1073
rect 835 -1085 841 -1080
rect 987 -1159 993 -1153
rect 835 -1167 841 -1162
rect 632 -1310 639 -1303
rect 926 -1318 936 -1310
rect 835 -1325 841 -1319
rect 1061 -1235 1067 -1229
rect 1077 -1241 1083 -1236
rect 1077 -1317 1083 -1311
<< m123contact >>
rect 887 -863 897 -855
rect 773 -1131 783 -1125
rect 889 -1249 896 -1243
rect 879 -1256 885 -1251
rect 869 -1263 875 -1257
rect 860 -1270 865 -1265
<< metal3 >>
rect 78 -1091 85 -1057
rect 89 -1091 96 -963
rect 101 -1091 108 -871
rect 112 -1091 119 -779
rect 71 -1096 273 -1091
rect 78 -1369 85 -1096
rect 89 -1294 96 -1096
rect 101 -1219 108 -1096
rect 112 -1144 119 -1096
rect 112 -1151 225 -1144
rect 101 -1226 224 -1219
rect 89 -1301 224 -1294
rect 337 -1319 343 -761
rect 464 -814 866 -809
rect 464 -815 635 -814
rect 819 -815 866 -814
rect 349 -1333 354 -1142
rect 358 -1303 363 -853
rect 464 -879 471 -815
rect 367 -1288 372 -1215
rect 386 -1359 391 -884
rect 400 -1032 405 -893
rect 464 -935 471 -885
rect 400 -1033 406 -1032
rect 405 -1038 406 -1033
rect 400 -1347 406 -1038
rect 410 -1091 414 -991
rect 410 -1329 415 -1096
rect 464 -1156 471 -942
rect 486 -827 619 -821
rect 486 -888 492 -827
rect 475 -1020 482 -1005
rect 475 -1076 482 -1027
rect 486 -1069 492 -893
rect 594 -916 603 -888
rect 620 -903 626 -828
rect 498 -923 603 -916
rect 498 -975 505 -923
rect 498 -1062 505 -994
rect 620 -1012 626 -920
rect 632 -1019 639 -926
rect 801 -960 806 -905
rect 669 -966 806 -960
rect 475 -1148 482 -1083
rect 604 -1106 610 -1070
rect 502 -1112 610 -1106
rect 632 -1105 639 -1025
rect 502 -1235 508 -1112
rect 604 -1188 610 -1156
rect 512 -1194 610 -1188
rect 512 -1228 518 -1194
rect 632 -1303 639 -1111
rect 669 -1188 675 -966
rect 706 -975 751 -972
rect 691 -977 751 -975
rect 817 -976 824 -886
rect 691 -981 712 -977
rect 800 -1053 805 -1010
rect 682 -1058 805 -1053
rect 682 -1182 687 -1058
rect 705 -1071 710 -1065
rect 817 -1073 824 -983
rect 773 -1132 781 -1131
rect 691 -1137 781 -1132
rect 691 -1175 696 -1137
rect 817 -1310 824 -1079
rect 835 -986 841 -893
rect 859 -962 866 -815
rect 1011 -924 1016 -864
rect 870 -930 1016 -924
rect 835 -1080 841 -991
rect 870 -1013 876 -930
rect 835 -1162 841 -1085
rect 835 -1319 841 -1167
rect 860 -1019 876 -1013
rect 860 -1265 865 -1019
rect 999 -1025 1004 -970
rect 870 -1030 1004 -1025
rect 870 -1257 875 -1030
rect 999 -1031 1004 -1030
rect 993 -1111 999 -1072
rect 879 -1116 999 -1111
rect 879 -1251 884 -1116
rect 905 -1124 955 -1120
rect 987 -1199 993 -1159
rect 889 -1206 993 -1199
rect 889 -1243 895 -1206
rect 860 -1318 926 -1311
rect 860 -1329 868 -1318
rect 1061 -1322 1067 -1235
rect 1077 -1311 1083 -1241
rect 410 -1336 868 -1329
rect 875 -1328 1067 -1322
rect 875 -1342 881 -1328
rect 578 -1347 881 -1342
rect 400 -1348 881 -1347
rect 400 -1354 585 -1348
rect 78 -1376 224 -1369
rect 78 -1377 231 -1376
<< m4contact >>
rect 336 -748 343 -741
rect 172 -769 179 -762
rect 159 -861 166 -854
rect 146 -953 153 -946
rect 134 -1046 141 -1039
rect 225 -1140 230 -1135
rect 224 -1214 229 -1209
rect 224 -1289 229 -1284
rect 358 -787 367 -779
rect 444 -884 450 -879
rect 509 -991 514 -986
rect 658 -988 665 -982
rect 607 -1239 613 -1234
rect 784 -1186 791 -1181
rect 1080 -937 1086 -931
rect 1080 -948 1087 -941
rect 1020 -1035 1028 -1027
rect 1081 -1043 1086 -1038
rect 1213 -1085 1220 -1079
rect 996 -1254 1001 -1249
rect 996 -1353 1001 -1346
rect 224 -1364 229 -1359
rect 607 -1366 613 -1360
rect 659 -1369 665 -1362
rect 785 -1364 792 -1355
rect 785 -1383 793 -1375
<< metal4 >>
rect -94 -1329 -80 -531
rect 343 -748 1084 -741
rect 134 -1359 141 -1046
rect 146 -1284 153 -953
rect 159 -1209 166 -861
rect 172 -1135 179 -769
rect 367 -780 471 -779
rect 367 -787 1028 -780
rect 442 -788 694 -787
rect 444 -929 450 -884
rect 444 -934 514 -929
rect 509 -986 514 -934
rect 658 -982 665 -981
rect 658 -989 665 -988
rect 172 -1140 225 -1135
rect 159 -1214 224 -1209
rect 146 -1289 224 -1284
rect 134 -1364 224 -1359
rect 607 -1360 613 -1239
rect 659 -1362 665 -989
rect 1020 -1027 1028 -787
rect 1080 -931 1084 -748
rect 1080 -984 1085 -948
rect 1080 -987 1257 -984
rect 1081 -1081 1085 -1043
rect 1081 -1085 1213 -1081
rect 785 -1181 791 -1180
rect 785 -1355 791 -1186
rect 996 -1346 1001 -1254
rect 1250 -1350 1257 -987
rect 1065 -1358 1257 -1350
rect 785 -1419 793 -1383
rect 1065 -1419 1073 -1358
rect 785 -1426 1073 -1419
<< m5contact >>
rect 579 -912 585 -905
rect 1001 -910 1009 -903
rect 707 -944 714 -938
rect 570 -1017 576 -1010
rect 594 -1100 600 -1093
rect 229 -1168 237 -1160
rect 585 -1183 591 -1176
rect 228 -1243 236 -1235
rect 519 -1277 526 -1270
rect 582 -1275 588 -1268
rect 228 -1318 236 -1310
rect 989 -1009 997 -1002
rect 1089 -978 1097 -970
rect 707 -1041 714 -1035
rect 1089 -1076 1097 -1068
rect 980 -1102 988 -1095
rect 706 -1129 713 -1123
rect 1089 -1176 1097 -1168
rect 967 -1186 974 -1180
rect 704 -1228 711 -1222
rect 904 -1305 911 -1299
rect 984 -1304 991 -1298
rect 1089 -1274 1097 -1266
rect 996 -1377 1001 -1370
rect 228 -1393 236 -1385
rect 292 -1393 298 -1386
<< metal5 >>
rect 1260 -633 1315 -628
rect -362 -928 -335 -727
rect 186 -810 232 -802
rect 186 -894 195 -810
rect 186 -902 222 -894
rect -362 -934 -297 -928
rect -362 -938 -335 -934
rect -362 -947 -101 -938
rect -362 -1118 -335 -947
rect 186 -986 195 -902
rect 579 -927 585 -912
rect 579 -933 602 -927
rect 597 -939 602 -933
rect 597 -944 707 -939
rect 186 -994 226 -986
rect 186 -1079 195 -994
rect 217 -995 226 -994
rect 597 -996 602 -944
rect 1001 -955 1006 -910
rect 1260 -930 1269 -633
rect 1472 -784 1493 -607
rect 1379 -791 1493 -784
rect 1274 -824 1318 -817
rect 1001 -960 1016 -955
rect 570 -1002 656 -996
rect 570 -1010 576 -1002
rect 649 -1036 656 -1002
rect 1011 -1004 1016 -960
rect 997 -1009 1016 -1004
rect 649 -1041 707 -1036
rect 186 -1087 218 -1079
rect 649 -1080 656 -1041
rect 596 -1086 656 -1080
rect -362 -1125 -303 -1118
rect -362 -1129 -335 -1125
rect -362 -1138 -101 -1129
rect -362 -1313 -335 -1138
rect 186 -1160 195 -1087
rect 596 -1093 602 -1086
rect 600 -1100 602 -1093
rect 547 -1117 588 -1116
rect 547 -1122 584 -1117
rect 596 -1136 602 -1100
rect 1011 -1096 1016 -1009
rect 988 -1102 1016 -1096
rect 656 -1129 706 -1124
rect 656 -1136 660 -1129
rect 596 -1142 660 -1136
rect 186 -1168 229 -1160
rect 186 -1235 195 -1168
rect 596 -1178 602 -1142
rect 591 -1183 602 -1178
rect 186 -1243 228 -1235
rect 186 -1310 195 -1243
rect 596 -1270 602 -1183
rect 1011 -1182 1016 -1102
rect 974 -1186 1016 -1182
rect 970 -1187 1016 -1186
rect 704 -1270 710 -1228
rect 588 -1275 710 -1270
rect -362 -1318 -303 -1313
rect -119 -1318 -96 -1310
rect 186 -1318 228 -1310
rect -362 -1322 -335 -1318
rect -119 -1322 -109 -1318
rect -362 -1329 -109 -1322
rect -362 -1509 -335 -1329
rect -194 -1351 -137 -1342
rect 186 -1385 195 -1318
rect 186 -1393 228 -1385
rect 519 -1386 525 -1277
rect 704 -1300 710 -1275
rect 704 -1304 904 -1300
rect 1011 -1299 1016 -1187
rect 1045 -978 1089 -970
rect 1045 -1068 1056 -978
rect 1274 -1029 1283 -824
rect 1472 -974 1493 -791
rect 1389 -980 1493 -974
rect 1045 -1076 1089 -1068
rect 1045 -1168 1056 -1076
rect 1472 -1162 1493 -980
rect 1045 -1176 1089 -1168
rect 1388 -1169 1493 -1162
rect 1045 -1266 1056 -1176
rect 1045 -1274 1089 -1266
rect 991 -1304 1016 -1299
rect 1472 -1323 1493 -1169
rect 1408 -1330 1493 -1323
rect 1001 -1377 1318 -1370
rect 1313 -1385 1318 -1377
rect 298 -1393 525 -1386
rect -304 -1509 -297 -1498
rect -99 -1509 -93 -1495
rect 186 -1509 195 -1393
rect -362 -1510 195 -1509
rect -362 -1518 196 -1510
rect 174 -1563 196 -1518
rect 1384 -1563 1391 -1542
rect 1472 -1562 1493 -1330
rect 1472 -1563 1492 -1562
rect 172 -1591 1492 -1563
<< m6contact >>
rect 218 -731 226 -723
rect 218 -823 226 -815
rect 907 -834 915 -826
rect 578 -853 586 -845
rect 706 -875 714 -867
rect 218 -915 226 -907
rect 906 -940 914 -932
rect 568 -954 576 -946
rect 706 -980 714 -972
rect 218 -1008 226 -1000
rect 593 -1039 601 -1031
rect 906 -1041 914 -1033
rect 705 -1071 713 -1063
rect 227 -1111 236 -1102
rect 584 -1125 592 -1117
rect 904 -1128 912 -1120
rect 226 -1186 235 -1177
rect 703 -1153 711 -1145
rect 584 -1205 592 -1197
rect 226 -1261 235 -1252
rect 903 -1222 911 -1214
rect 226 -1336 235 -1327
<< metal6 >>
rect -266 -948 -250 -540
rect 1067 -617 1275 -603
rect -152 -731 218 -723
rect 226 -727 251 -723
rect 226 -728 261 -727
rect -152 -774 -137 -731
rect -184 -780 -137 -774
rect -152 -793 -137 -780
rect -152 -800 -96 -793
rect -266 -1140 -255 -953
rect -152 -963 -137 -800
rect 202 -815 210 -731
rect 224 -815 258 -814
rect 202 -823 218 -815
rect 226 -819 258 -815
rect 226 -820 263 -819
rect 202 -906 210 -823
rect 908 -826 937 -825
rect 899 -834 907 -826
rect 915 -831 937 -826
rect 1067 -826 1076 -617
rect 1006 -833 1076 -826
rect 1001 -834 1076 -833
rect 899 -845 905 -834
rect 1001 -835 1019 -834
rect 558 -851 578 -846
rect 586 -850 905 -845
rect 202 -907 259 -906
rect 202 -915 218 -907
rect 226 -911 259 -907
rect -186 -971 -137 -963
rect -152 -976 -137 -971
rect -152 -982 2 -976
rect -263 -1331 -256 -1147
rect -152 -1158 -137 -982
rect 202 -999 210 -915
rect 552 -953 568 -947
rect 607 -947 612 -850
rect 691 -868 696 -850
rect 691 -875 706 -868
rect 714 -873 742 -867
rect 576 -952 612 -947
rect 202 -1000 256 -999
rect 202 -1008 218 -1000
rect 226 -1004 256 -1000
rect 202 -1102 210 -1008
rect 607 -1031 612 -952
rect 691 -972 697 -875
rect 900 -932 905 -850
rect 1065 -891 1076 -834
rect 1267 -637 1275 -617
rect 1356 -620 1362 -533
rect 1267 -645 1326 -637
rect 1267 -826 1275 -645
rect 1356 -810 1362 -626
rect 1267 -834 1331 -826
rect 1267 -844 1275 -834
rect 1065 -896 1095 -891
rect 1065 -900 1098 -896
rect 900 -940 906 -932
rect 914 -937 939 -932
rect 691 -980 706 -972
rect 714 -977 743 -972
rect 691 -981 714 -980
rect 555 -1037 593 -1031
rect 601 -1039 612 -1031
rect 606 -1054 612 -1039
rect 606 -1059 619 -1054
rect 224 -1102 262 -1101
rect 202 -1111 227 -1102
rect 236 -1107 262 -1102
rect -187 -1159 -137 -1158
rect -187 -1165 1 -1159
rect -187 -1166 -137 -1165
rect -152 -1339 -137 -1166
rect 202 -1177 210 -1111
rect 550 -1117 588 -1116
rect 614 -1117 619 -1059
rect 691 -1063 697 -981
rect 900 -1033 905 -940
rect 1065 -989 1076 -900
rect 1065 -994 1090 -989
rect 1312 -994 1341 -988
rect 1065 -998 1097 -994
rect 911 -1033 949 -1032
rect 900 -1041 906 -1033
rect 914 -1038 949 -1033
rect 691 -1071 705 -1063
rect 713 -1068 735 -1063
rect 550 -1122 584 -1117
rect 592 -1122 619 -1117
rect 202 -1186 226 -1177
rect 235 -1182 264 -1177
rect 202 -1252 210 -1186
rect 614 -1197 619 -1122
rect 691 -1145 697 -1071
rect 900 -1118 905 -1041
rect 1065 -1089 1076 -998
rect 1333 -1017 1341 -994
rect 1356 -999 1362 -815
rect 1335 -1022 1341 -1017
rect 1226 -1080 1245 -1077
rect 1232 -1089 1245 -1080
rect 1065 -1094 1095 -1089
rect 1226 -1094 1245 -1089
rect 1065 -1098 1101 -1094
rect 900 -1120 943 -1118
rect 900 -1128 904 -1120
rect 912 -1124 943 -1120
rect 691 -1153 703 -1145
rect 711 -1150 730 -1145
rect 555 -1203 584 -1197
rect 592 -1203 619 -1197
rect 900 -1213 906 -1128
rect 1014 -1137 1030 -1136
rect 1014 -1146 1023 -1137
rect 1014 -1149 1026 -1146
rect 900 -1214 959 -1213
rect 900 -1222 903 -1214
rect 911 -1218 959 -1214
rect 231 -1252 263 -1251
rect 202 -1261 226 -1252
rect 235 -1257 263 -1252
rect 268 -1257 269 -1251
rect 202 -1327 210 -1261
rect 234 -1327 263 -1326
rect 202 -1336 226 -1327
rect 235 -1332 263 -1327
rect -152 -1340 5 -1339
rect -152 -1342 2 -1340
rect -189 -1346 2 -1342
rect -189 -1350 -137 -1346
rect -194 -1351 -137 -1350
rect 1014 -1359 1023 -1149
rect 1065 -1187 1076 -1098
rect 1065 -1192 1092 -1187
rect 1065 -1196 1099 -1192
rect 1235 -1207 1241 -1094
rect 1356 -1188 1362 -1005
rect 1235 -1212 1329 -1207
rect 1046 -1337 1062 -1334
rect 1235 -1337 1241 -1212
rect 1046 -1344 1298 -1337
rect 1061 -1346 1298 -1344
rect 1061 -1351 1062 -1346
rect 1014 -1387 1024 -1359
rect 1286 -1395 1298 -1346
rect 1356 -1376 1362 -1194
rect 1286 -1400 1327 -1395
<< pad >>
rect -269 -540 -247 -532
rect -93 -538 -74 -532
rect 1354 -533 1364 -527
rect -305 -934 -296 -927
rect 251 -727 262 -722
rect -95 -768 -79 -760
rect 172 -769 181 -762
rect -197 -780 -184 -774
rect -100 -779 -76 -773
rect 112 -780 120 -772
rect -96 -800 -88 -793
rect -267 -953 -248 -948
rect -304 -1125 -297 -1118
rect 218 -778 226 -771
rect 224 -809 234 -799
rect 258 -819 264 -814
rect 24 -862 31 -852
rect 159 -861 166 -854
rect 618 -830 628 -819
rect 937 -834 944 -822
rect 999 -833 1006 -825
rect 356 -857 368 -846
rect 552 -852 558 -844
rect 384 -885 393 -878
rect 462 -885 471 -877
rect 476 -882 486 -876
rect 593 -886 602 -879
rect 218 -901 224 -894
rect 400 -896 407 -887
rect 485 -894 493 -889
rect 259 -913 266 -906
rect 579 -912 585 -906
rect -108 -947 -101 -939
rect 50 -955 61 -944
rect 146 -953 153 -946
rect -95 -963 -80 -957
rect -197 -971 -186 -963
rect -184 -1028 -177 -1023
rect -268 -1147 -252 -1140
rect -304 -1318 -298 -1313
rect 2 -983 10 -975
rect 462 -942 473 -935
rect 546 -954 552 -946
rect 742 -875 750 -866
rect 620 -909 628 -901
rect 638 -904 646 -897
rect 620 -920 627 -914
rect 634 -927 643 -921
rect 497 -981 506 -973
rect 222 -993 228 -986
rect 407 -992 417 -985
rect 497 -994 506 -987
rect 571 -990 582 -981
rect 256 -1005 266 -998
rect 422 -1008 432 -998
rect 476 -1005 484 -998
rect 54 -1046 65 -1036
rect 133 -1047 141 -1039
rect 569 -1016 579 -1010
rect 473 -1028 481 -1023
rect 399 -1039 406 -1032
rect 549 -1038 555 -1030
rect 815 -888 825 -877
rect 846 -878 854 -870
rect 834 -895 842 -887
rect 799 -907 809 -898
rect 1009 -866 1017 -857
rect 1354 -626 1363 -620
rect 1310 -631 1315 -626
rect 1326 -646 1334 -635
rect 1379 -791 1388 -784
rect 1354 -815 1364 -810
rect 1312 -821 1318 -816
rect 1331 -836 1336 -826
rect 1095 -896 1103 -890
rect 999 -910 1010 -901
rect 705 -946 717 -937
rect 939 -939 946 -931
rect 862 -969 868 -961
rect 743 -978 752 -970
rect 618 -1019 629 -1012
rect 634 -1028 642 -1020
rect 618 -1049 627 -1041
rect 504 -1066 510 -1060
rect 489 -1074 499 -1069
rect 218 -1087 227 -1079
rect 476 -1085 486 -1080
rect 409 -1097 415 -1089
rect 592 -1100 600 -1092
rect 262 -1109 269 -1101
rect -108 -1138 -101 -1130
rect -95 -1145 -80 -1140
rect -195 -1166 -187 -1158
rect 1 -1166 11 -1157
rect -185 -1223 -176 -1214
rect -264 -1336 -255 -1331
rect 544 -1122 550 -1116
rect 814 -985 827 -975
rect 847 -977 856 -970
rect 834 -992 843 -985
rect 798 -1011 807 -1003
rect 997 -972 1006 -964
rect 1082 -937 1089 -931
rect 1262 -932 1270 -923
rect 1081 -949 1088 -942
rect 1090 -994 1104 -989
rect 1304 -994 1312 -988
rect 987 -1011 997 -1001
rect 705 -1041 716 -1034
rect 949 -1039 956 -1032
rect 1019 -1037 1028 -1026
rect 735 -1071 743 -1061
rect 805 -1068 814 -1061
rect 643 -1102 651 -1095
rect 627 -1111 638 -1105
rect 225 -1151 232 -1144
rect 478 -1152 488 -1146
rect 598 -1157 607 -1149
rect 228 -1168 237 -1160
rect 462 -1164 472 -1157
rect 264 -1184 271 -1176
rect 583 -1182 591 -1175
rect 815 -1080 824 -1073
rect 833 -1086 842 -1079
rect 992 -1073 1000 -1065
rect 1384 -981 1392 -974
rect 1353 -1005 1364 -999
rect 1331 -1022 1335 -1017
rect 1274 -1029 1282 -1022
rect 1081 -1046 1097 -1037
rect 1224 -1089 1232 -1080
rect 1095 -1094 1106 -1089
rect 979 -1104 990 -1094
rect 705 -1131 715 -1122
rect 943 -1125 955 -1118
rect 730 -1153 740 -1144
rect 833 -1170 845 -1160
rect 543 -1205 555 -1197
rect 1023 -1146 1031 -1137
rect 986 -1160 994 -1151
rect 967 -1189 975 -1179
rect 513 -1231 521 -1224
rect 703 -1229 711 -1221
rect 959 -1219 965 -1209
rect 228 -1244 237 -1235
rect 499 -1242 511 -1236
rect 263 -1257 268 -1249
rect 498 -1253 510 -1247
rect 994 -1255 1002 -1248
rect -104 -1318 -97 -1310
rect -95 -1330 -80 -1323
rect 518 -1276 528 -1270
rect 580 -1276 588 -1268
rect 641 -1284 650 -1277
rect 226 -1316 238 -1310
rect 629 -1313 641 -1301
rect 813 -1311 821 -1306
rect 832 -1325 842 -1317
rect 925 -1319 938 -1309
rect 263 -1333 268 -1326
rect -195 -1350 -189 -1341
rect 2 -1347 11 -1340
rect 994 -1354 1003 -1345
rect 780 -1383 801 -1355
rect 1089 -1144 1096 -1137
rect 1092 -1192 1104 -1186
rect 1379 -1170 1392 -1161
rect 1355 -1194 1363 -1188
rect 1329 -1213 1334 -1205
rect 1045 -1357 1061 -1344
rect 227 -1394 238 -1385
rect 290 -1394 301 -1385
rect 1011 -1394 1025 -1387
rect 1405 -1330 1413 -1323
rect 1311 -1385 1319 -1380
rect 1355 -1383 1363 -1376
rect -182 -1405 -175 -1399
rect 1327 -1400 1332 -1394
rect -303 -1504 -297 -1498
rect -99 -1500 -93 -1495
rect 1384 -1549 1392 -1540
<< labels >>
rlabel metal1 322 -945 336 -940 1 p1
rlabel metal1 322 -1038 336 -1033 1 p0
rlabel metal1 290 -1139 308 -1135 1 g3
rlabel metal1 288 -1214 315 -1210 1 g2
rlabel metal1 289 -1289 316 -1285 1 g1
rlabel metal1 289 -1364 314 -1360 1 g0
rlabel metal1 162 -767 165 -764 1 A_3
rlabel metal1 105 -776 107 -774 1 B_3
rlabel metal1 90 -867 92 -866 1 B_2
rlabel metal1 99 -858 103 -856 1 A_2
rlabel metal1 90 -950 93 -950 1 A_1
rlabel metal1 83 -959 85 -958 1 B_1
rlabel metal1 81 -1045 84 -1041 1 A_0
rlabel metal1 67 -1053 69 -1052 1 B_0
rlabel space 322 -854 337 -848 1 p2
rlabel space 321 -762 343 -756 1 p3
rlabel metal1 608 -1373 611 -1371 1 CARRY_2
rlabel metal1 660 -1378 663 -1374 1 CARRY_1
rlabel metal1 786 -1373 787 -1372 1 CARRY_3
rlabel metal6 213 -731 226 -723 5 vdd
rlabel metal3 71 -1096 77 -1091 1 C_0
rlabel metal1 -109 -786 -107 -785 1 b3
rlabel metal1 -304 -767 -302 -765 1 a3
rlabel metal1 -306 -957 -305 -956 1 a2
rlabel metal1 -108 -969 -106 -967 1 b2
rlabel metal1 -104 -1152 -102 -1150 1 b1
rlabel metal1 -305 -1152 -304 -1150 1 a1
rlabel metal1 -306 -1336 -305 -1334 1 a0
rlabel metal1 -101 -1333 -100 -1332 1 b0
rlabel space -294 -504 -154 -473 1 clk
rlabel pad 218 -901 224 -894 1 gnd
rlabel metal1 1448 -699 1452 -697 1 sum3
rlabel metal1 1454 -1456 1460 -1453 1 CARRY_4
rlabel metal1 1448 -1268 1455 -1266 1 sum0
rlabel metal1 1455 -1079 1458 -1077 1 sum1
rlabel metal1 1454 -889 1456 -887 1 sum2
<< end >>
